module uart_top(wb_clk_i, wb_rst_i, wb_adr_i, wb_dat_i, wb_dat_o, wb_we_i,
	wb_stb_i, wb_cyc_i, wb_ack_o, wb_sel_i, int_o, stx_pad_o, srx_pad_i,
	rts_pad_o, cts_pad_i, dtr_pad_o, dsr_pad_i, ri_pad_i, dcd_pad_i);
	parameter		uart_data_width	= 32;
	parameter		uart_addr_width	= 5;
	input			wb_clk_i;
	input			wb_rst_i;
	input			wb_we_i;
	input			wb_stb_i;
	input			wb_cyc_i;
	output			wb_ack_o;
	output			int_o;
	input			srx_pad_i;
	input			cts_pad_i;
	input			dsr_pad_i;
	input			ri_pad_i;
	input			dcd_pad_i;
	output			stx_pad_o;
	output			rts_pad_o;
	output			dtr_pad_o;
	input	[(uart_addr_width - 1):0]
				wb_adr_i;
	input	[(uart_data_width - 1):0]
				wb_dat_i;
	output	[(uart_data_width - 1):0]
				wb_dat_o;

	wire	[7:0]		wb_dat8_i;
	wire	[7:0]		wb_dat8_o;
	wire	[31:0]		wb_dat32_o;
	input	[3:0]		wb_sel_i;
	wire	[(uart_addr_width - 1):0]
				wb_adr_int;
	wire			we_o;
	wire			re_o;
	wire	[3:0]		ier;
	wire	[3:0]		iir;
	wire	[1:0]		fcr;
	wire	[4:0]		mcr;
	wire	[7:0]		lcr;
	wire	[7:0]		msr;
	wire	[7:0]		lsr;
	wire	[(8 - 1):0]	rf_count;
	wire	[(8 - 1):0]	tf_count;
	wire	[2:0]		tstate;
	wire	[3:0]		rstate;
	uart_wb wb_interface(
		.clk				(wb_clk_i), 
		.wb_rst_i			(wb_rst_i), 
		.wb_dat_i			(wb_dat_i), 
		.wb_dat_o			(wb_dat_o), 
		.wb_dat8_i			(wb_dat8_i), 
		.wb_dat8_o			(wb_dat8_o), 
		.wb_sel_i			(wb_sel_i), 
		.wb_dat32_o			(wb_dat32_o), 
		.wb_we_i			(wb_we_i), 
		.wb_stb_i			(wb_stb_i), 
		.wb_cyc_i			(wb_cyc_i), 
		.wb_ack_o			(wb_ack_o), 
		.wb_adr_i			(wb_adr_i), 
		.wb_adr_int			(wb_adr_int), 
		.we_o				(we_o), 
		.re_o				(re_o));
	uart_regs regs(
		.clk				(wb_clk_i), 
		.wb_rst_i			(wb_rst_i), 
		.wb_addr_i			(wb_adr_int), 
		.wb_dat_i			(wb_dat8_i), 
		.wb_dat_o			(wb_dat8_o), 
		.wb_we_i			(we_o), 
		.wb_re_i			(re_o), 
		.modem_inputs			({cts_pad_i, dsr_pad_i,
		ri_pad_i, dcd_pad_i}), 
		.stx_pad_o			(stx_pad_o), 
		.srx_pad_i			(srx_pad_i), 
		.ier				(ier), 
		.iir				(iir), 
		.fcr				(fcr), 
		.mcr				(mcr), 
		.lcr				(lcr), 
		.msr				(msr), 
		.lsr				(lsr), 
		.rf_count			(rf_count), 
		.tf_count			(tf_count), 
		.tstate				(tstate), 
		.rstate				(rstate), 
		.rts_pad_o			(rts_pad_o), 
		.dtr_pad_o			(dtr_pad_o), 
		.int_o				(int_o));
	uart_debug_if dbg(
		.wb_dat32_o			(wb_dat32_o[31:0]), 
		.wb_adr_i			(wb_adr_int[(5 - 1):0]), 
		.ier				(ier[3:0]), 
		.iir				(iir[3:0]), 
		.fcr				(fcr[1:0]), 
		.mcr				(mcr[4:0]), 
		.lcr				(lcr[7:0]), 
		.msr				(msr[7:0]), 
		.lsr				(lsr[7:0]), 
		.rf_count			(rf_count[(8 - 1):0]), 
		.tf_count			(tf_count[(8 - 1):0]), 
		.tstate				(tstate[2:0]), 
		.rstate				(rstate[3:0]));

	initial begin
	  $display(
		  "(%m) UART INFO: Data bus width is 32. Debug Interface present.\n"
		  );
	  $display("(%m) UART INFO: Doesn't have baudrate output\n");
	end
endmodule

`protected
g<HZ8e25S&O+:35C1U6ae+HdE6CBL<A@WV9#7+JNg5R_b2C[Dc+g4)T+(0B8_gDW
bT71>MYTWKA@U&/4/V9QN-K,B3G)F=M0CTEeJXK#ECd=4S+BN\TMP2P);C4;F&\C
#?Z2dBPVB2#^)eQ+9P;a1aQ862;7)1+;<g2D(>4YN3E?##9.E_\AW/P<:AG?_B_C
J2WT<]T[B@68=/WX6R01GgMP5WI^-2J:CJ66?V;[C:-Ka8B2__FALX@b;,D;:..]
1]_ATd#8,Ra7F<A=+b]F\5/(2RKg46DR+cc26e3,OQF^H?L[Q^?[Ug>1ZVBIV8;.
Yg=@e6E+2+[<YR2@TIa&&]K.@GVOe;-RYGa/#&(D@G><IOIPDO+6IC[J2@PZJU;e
QADg-RT?Z[eF8B1Df3F5I?MQSgHYM#bSRY,B>:Q710+fOa7.ce/AYPNNfRX-3:/[
c7,RYbJaCS:CFecXYRK=Me1)H5CJ+M(4,6OR1<_:VU],];57Q#^4G@Yg2XGScF+P
cbS^=dQeP.WdNNZ^S\&R@9M>AXLL1>P6:(;]U_PW3RgXHETOLUdSfgZTLF_PJAYR
CZ<OGX+C5WHNTg>Q0046c;>CV1WJ&B)3?+F7B?-AFE.X,MUGdRaaeKG/d10?g>F4
Z<g/eCL5J2^]:TMVM9R>A,E[gQNR[,C_CZ/QC#ge\8>.=I1MYSN0d[072Z.W,+\9
(26(D17gR^d[MVS^QYb?1UQQV+R\cM9UQFb[Q[V(RO<S-DA.)gb/9HPBHV-D20#C
I1QHBG4F1dT6d<aV/FePJ=:HZ4E24RPQ33CD(DfeO(/>)W@fD\:8T(8SHES@BD4O
cC?>aFDHO9<&_.@]&EaSY(AU#Ud\)S.=JHCdbY]#F#_ROcO+&e8E8E3QQ\<#/1JA
2>XI6@)Eg4SKUVLG/Ua=E-PWc])_c?OI^\.^7,4[<):g5Y9L#YU5#N\,CZg7NeHd
(S]OG:O[0H\H[Id?^Of8UM-bP&&1X[Qgf2MU3&H=YRT5<XCN69QL8_ZYL;G/1R]K
:GK@;GV^e)bf3&VNa>]?-E3eN5N5a^IJ#_[2Yc+V2X?gXE+bZQ^JIXd;19[(,QAb
+<JZ8SG6PVPF>RIJ,\G\AOT6)=<GK(dXIe(D(R8F3aATK]ZMb5cV,NKV=a6GVEJP
-7_5TPb3#1/-AbN#=Z_0OERf75=SU?\eE?QHT1[g^9b5eNH@:=NHcQNU6R]Y&RB@
AUFGIZ^V2W>#>=^_=(&<gEe^2[3&G:C)IY;(_1g]bHFN1^e&B7K=3ZdYR]P[\e]\
JdOHd)]JB21Y+WW,=;aU\YOMa]Vf+SF(eD0[,1&2FF.bVR^Q=ZaJWd/RFWMKc[Q1
]a_[(KA3=]&90BEZ2eEQ5OZ?<R7+9_1BGW+K7U>EF;R.):gGgTLYZ322)RQ?=K2Q
A4N7c_\VMOZ0Vc05@M9/e_8?S^a1EbDPK3TD95QfdZQ8U_,f8D/CBJY)0+fA]P#M
AK7C>QFLBJ7SedA>eg5V+S79<E^,L[+Jf1K10KM2<-G&-CB_4UQ@_37E1Ped@-/F
X&[cY>[75QK/(=6SY_A?X0_L?.G0VF)]E/YUT..Ue^]<.FG75,SE^K+-YQ<GR#/;
G:>@(AaIaD559?J21gK7?.B=[d&#7Z<68e,,ZcW/9dP_+ed)(VbX87d2,8^d\BGA
A-WY9;N0_COc:Y@=)&#4WVNg^T.NV.0F#bB[f>NK&S9:()()g\[(9QPQ_LCf>+#W
dC#<<U#HXU2HLN4AL[/LFe?)RZE43S.g=U3:DGS1E;#HP[AgNGGSA_fdaT_#(N;F
TS9&K)\7[G#]??f/AN9T787VbVC[\@PQ/PP>=<)4UD;V_>ITE?Q9a2a6=<?,7G61
?<@H&42/a]7G>W:3CW+P+f_=5K)F/I@@RN)9Z2gc43REgRE,cJ](2M@aR#C#a9]B
+^^GC@fb:\999>^O,7@[TFY70X=N(I23AC]-edf<,+6d3.ga<\CM4)PT[gQ53dQ]
K.&_VM8/MK\:ec0f9UAe-45LZIDbMAGIDL:GJ<L9^Gc/YbR]9ICUC@7K@69(:&]D
7(4eJO#06K-+FQ=&8;gI@T&@H^(=dMD1B)R&UL7Q5QAdD?MX=NY6;=?]&O8S#>D&
=7+Jf_YbZ<;&IS6:+UV]>Z?#_eKVGF]GaE8E-b0PQJ8(581C)]_dU/>XK(-ELBWa
ZY@Oa:DAED-?aK][7N8A4d<gY5CX>5QfOUA+(,6(P3.VCVdJ&\8T@U]410Q83Y6A
NLG#(&9JWGZ;IO3IG;-dJR906]LT)agP&RG[V5TR8T7_11V^WDU9aVYZ=0<J5_BL
/4_6F/+ST>7AJA69X.a.e@:_>8B-Z3I->H77ffbHHaFA#3[N-Y,\4;C=R0K@1A\a
GbWSeLf-KQ(W@H_Y2=0,BbIJPG5&ON/aV;,YX@N4>8;7E&C15eL^SDa(68RCX,)X
6S>TYe&>UAH#9_O^,YH5T8-.>]TA9g1JGO.@Q[^9-]dLO:[[[5PdGYNONOSbb;&C
10?fXH:1eWGPW2HB#L)]<TESO4ZG/K-WICE^U@8Q&?E-OS97gE2PK-&?(>C(_1O@
)6(PSD^2b2eYe(8LXIG?-N[W0II94.cP-7-a7FaE-[9W,S.I^5S-2RX\RB]+&\1R
d;>CRU-XN\#WWRX]dK=)AA5GGDCYKPWSH6f_U;]ad-7K4[b03++A&?G1,Ub?]58?
/&O7O6?T<N9RLRFSRI86H/]A(ZX:L1\<aH]3UBGOBgb\QWH/^FS>eZQZR[W299/8
>#gX;O;6b@EAMN2^\/0#dNcRYTBX)d,[VU1g4?=<:ES#5.dVId6O&A>+QLZ;09I<
4ee13S[OSf)?[&08RELC7KEG<EB89@,_5J)(g(]b0Xg<=Q.#2a?ZQdY?WPNM8I+3
R[LeA[:+N6@M\,SHSgY]7>bQ/UL+0C:>)b\<04PKCD^gXK)H##H1PR0>>-K4J>?,
.SI7-O)K,V)T.U1SHW8Jc+PD.S-8GDH1AaTP(c21@CUDQAHF&[#T?,3_fS7<;OAL
8a;/N4_@[B9\XIDS]#3)[1>1R/ME,=6g#6JV33.HF<+gQIb2gX\[b+[(Z,AHL?fQ
c&\6O:>]9d:<P=4=?W70(NMH&EPd(\?JX@3fCfPEWC1M=TBJ^<X]2]T[cXe5HY0^
;8(e4<Z\SHcF6&=R[,5/WFdBcVL=fBBN766A0GC,=R,\Xfe9B9I]1+;AJY,b-1Q<
fF^a^]Y/0bI?L\Ve;4\A<<af/^aYDbXOL?GB/:=NR.M9MXZ.S/1+J)d^L_UFHV(T
)F@([U58Z5CYa86S?2;KC2X[&;g0KB,A)40C<+IN&)8]W\\9@#OAL.[Z_1(S2YUK
;EXMa7A=#\Y_WE\\A^+\Y;--C<>RaW&F:2_UEB-\eV018=e6D^,GG,F+9^W?5ZDc
=+-S6THBE3OI539XFQdF6GE83QJCRJ4#.M@,Ha)W:SATV&X;g-@KfaV,F[bPPL=T
5g0Z+@(VWCF]>S@9EBB-CEY+(US^ABdSPG0:<7>;_U/)R1EZGQO5]4/NW[QdH+=e
F2R)GO:b6N2PB4NRaQ/Cda\9H3^WD@\574J>BI^MQP&eNb(f7F@MdRBT?0-V5?Zf
@+?5RP_LK/\ZRW=4<NWcPDAQ?[F[G8@YY3(I6AfTP=dNT)61ZI?[6-//;K#NX:QS
IO<[EeXNe04g^=N=8>Z^X/^]?L9HPc-d>JeK:39EM:IC^GbcQP>BIX^;&D:PagcW
MR\a=8\;G->&[ZK+98-^A8=U#:RfQgY[IKbS>cg@YU4<Ig[,XaH;<f3HVM?^#&](
Zg+0FeU=G19++>g@2(G\fT/9dKS1g?2=;_=7-,?HQ+<OF^ec[DMH=TC61E[P,aQb
+6ceD3]LO7]9(0.@N454Z-f#gWD-GT3ee@/3KFO11^e&3F;>-D0d^1#::;9gcE4R
2-1.:N+H189Rb#D9F2\R]#_f/QZ-7E+>434H[-CR(QY>C?[C\AOBKL7XMS0S4_W3
Z_NMN[HCf=e-VA5BH5,\(/\0K[KVMCd?IVT^AYEC>CH^URPgUa>IHO@-/AD\LCfU
)>@DCPV4OQRQL48B6f5_^@?-E)8(Wc/-D64@@TO/,^gUPa0[X,g&\QTZW:e9QX<-
9D;4@<g,P(D;CMD/W:V=<U5gP3;>/]H8OBZZ;/9@/f&04U.>-RH5CeINF;82O^Yd
Q;Jg&.&>aSOEN\R:&R0(MDdL<ge:&3Y@S7)</_aKDJUSQ+6P8O,gYQ].U@@RT<NT
PHU\bVYN33<^_/dOPM_Q.Y)C6CE))4>/0#PZ[BGK+[@;3S=&)7@69@5G,?6S+ZE)
,FT(^:[XSS:4-+XGOR<0754+UeUPeWBg7Pa64^#9VX3^Wga+W@-F7Ua,1:@V/@F_
J_dQG9Vg#=,NMM.Z6PYW&=X<)\=5TLgE[W4-f:M6[b_<[,Y,2g]>80e9cD7YKbLa
9KYDX.B7R_;1P]:9I.YRX\TDafPd\McBJR6VHW;?XX;F#32B4_#:VC8b]]M_JLbY
?9=\f2ce)]S-X.9)KdYW9aC5RD?S\[7+&RA.OgYB)^:^TZPO<NX_/M[<(N:FG6XL
=@7ag@DID@<2Z++EbWN84<;La4,YSHR]N;G6D]ITUFK2IY>,e=MV2cW#8eAO\9fN
CFD91M@TFK9edPbaU(C-;G)T1G>P3Q0;?e++;7JSHZ3:A2E9fFI)K,B@&#VTf;g#
5gDg.F:3Add?2UggYW^R118_.0b\-?SD_<YHBG:.0-MBT>/FTIdI]0g-SDFX)Q+[
421JO54XQ6M5H3\07_Cf?IXcM&+6^THS^I#R#-/.\\,].]8)M,aQ-E,MAE2D\VY:
#;?K#8Sd-c;50#3aBdL3],[F7LD)RV>Q[E.L@<_S7OCGIgIb2WBUNOf<3LE,)-Y.
cX:A_Y/W:e.d)FJYE25)-C8\\OFUB>Z6gX>E8,/5<P@1#,dCKTJ/VZ5]ZQNc4UJF
:e69WJE,<BQMV2<^b4Q@)Bc\.;L/]bTU2_G?(b.:OV_G;6ee<//;E3B],dXZ^8Z)
ZJS-L]L)cId/J5<BbQ0U3E4eO++Q7S#@7HAa>Oa8-MdRC<N78#0?e;SY2_KTWSFW
)T@UWIe(:/-[)ET_4=U:;HaL4fDF/UCNPLM?SMWYV(c6NN7TbdGaTFSFBGF[7Q]K
A@OS^TGX.4a-X)[e-f\2RD^Z=aEX;B[@7)R=1L=RUB\5LHNCeSBEOW#8)a<(:Y4E
G1L(X+^e_Q;5@\OMQ&HKKU#_7X/\KF^D\+84=7&^H(#QF[T2?[JWTQ9;>K/T5R,L
2TVZ[-_<YgZ2\N.[7RfVe+T]+L.6437<[ZL4/<6S+bT^1+<H^G[BY;@@CVU=VE&g
e@-^5WgPefBIKa5d:BQUf2Q2A[a)eeB>LYM5c^U0+P2P:<\NgIB,CHSN.=X9>f@1
L^A=;#FDF=7]?AN?X<U\6&YZB6G#)>^&G30EA=a#d.6&f,NN.#9(]ENeS7ca?NQU
:2A0[aG@(dE21[\b6)<ed^5PWe0N:0H[)_>ZX59D:BS94RSb,::7S=-7Y8+YcU.I
0aM>(BJE1I4)_@V,27/NGDgc7GSOB;-,95Eg&DC7C0)EeHC#@1/f_L#Z>V.f68D0
5IT2XMe(^J6+=<:-^?g/QHO.7@P0YC1@deR6TX-P+4f1:ED:V#1CAO>e)RYBb>)E
X@/_X#;\9>=>D?=aH#K&5b;OC?aW,gAK(C-?Cd79KG7KU=VO^UMBBS=89O2H+IYa
bSddA46=CU1ADBe6fb.+1NP6<B^X^KF.X5G:_UL5\_B(3+/EIE,770>NK>]9F4P6
e7G#ScT42VIF6UB/]A/S1BDSgJ7+HAYJ=5B19a2Z1E_K8:g@HN0Cc?,;V4#HNBRa
CYB?9S9KGb#:I,X5:@I5E0g+B1U.T?T()\1G6-a^VEK+I2BddZddaUX@^aOOVeG-
K>c1M7cQeRLULW00#4e_3W<JT9=-.CJdW,NWaR@)/QG[1XHe]].A&&56d(HS&6W,
GJ<T.g]A7DfGA@F>VBdcB#C]E_ZQ);I&&P^#N:SL=\PYK<a9W@b.4geF;g0OC,UH
E&]gV>@X9B#.G0L?9^6SJba(/&,D/U(BD;Z)L<,eBf;#)Hb8QUC#BY1/dS>K</F@
0ITUf\Ua7eVE=?D:O]CSW=.,64ES):II.PJMRMJFD^MO9bP-\[7BW41H)@:JW^O6
0\e:C-e[JEUUVG=OY\OgU^b\dY0B?VWcZ>E<=F;;R2+2=VC#+1^NLeP-0@83:;TE
dG.SI?T+a2-Wg2NE>S64eOJ-E]b3WQCU,/>B]c<]K)KFRV&3X5VX&:)MbP+NUHc@
?c(Z8E@7OS>cSP4V0bG32Kg66gF;g#;F-,I6Jd\gB7)B#@B8UI-:=IY2f8GAg/V?
5#E5_GQL+-P7=2\.(H3I<S:g,-g;DYbS1>[8bGBSId=(N/c998N3^7\C1@34F.Jf
gIFaKM6aU8?IO6C_MCTOe<@++KHU#LKO8QRN,_e=(6[NcC1ILcE=I>P7D=,ffG>8
OJ39(,,e]@@],V_dBA+O5Y.FFTN+1f68fXd0)C.4VGMZX1E/>?.8A(W<&b,=B+TC
G5TebT+9->46;FdVM,5D]X4X#f2eO0Q<f+MNBb.:MK381,S6b,A4;MI>(#NPK6P_
B,@>Y#G6c<=E.LgK&,If:R>#5,AJ]f7X,g>[;F8eZ(C/fBF_CVaU5fKH3&E9b^]_
3+BXBb05[Y0eS]cR[BJ9UQ+a,8PeKWVdPfEgNC[AL&09AD;>\7N#)>FPd1/,KDc,
@)EHD/HddV7]^P6@>^O=RVBcJS3P7K/&Pbb\JCXMLY(Na#QFL06(N:e=-\a-@Y23
70c\Q;gN#^#67-+<6<Dd/N=JC7A-=L;5HP^7dd:J42C_S3H4GXFT?BD#A.ZA4gWQ
/;WQ#c1^Q^TO7->6J+G.)[2)_<WVRREBF7@>VX+PPAVFHME2#IGGDHJ?+3J^@7Vf
E.QIWCdHLY.4XdU;]5Ra>/.<+D;K:72?ga)-L>L+d_I3R8&WIC_@C@)/T8<I=CS=
@\cQ1Hg&d+BO5[OQc&@),9;+3=\L66?W2F&c<.)QYX:ZHCNI?g/7A8Gg55gZVL@g
LB1d&_;TaVGR\:4RI-)\NTYEJVQ[-cXNP&R2H,dX8TN(6<?]>P/BTQ<X:SRU21A5
?.NUY13BbJd.QK0YZ4QG[7SEB,gL:VRbQ1J)8>6/5^1Vd=R_63<U,D+1[PVYMWbC
WR?dda]#-6<NE>eZ?2MGF[I?e/IGHXfd:0R0:(J.)ZgRdVdeO5^48\U0Y5E6P6)[
&1N/\<_5BF:2N=;I+M,L(N(b8F=JFB/,)D948V;?75EWC6]N45d=TFGF^,eX-?>Q
C2WRa#NN?#HIaS^>J@MGBg@QCG=bg,9<7\Y7gNF8NVW8]XCF+B08M;]gF+Tc&(;Q
+2-3SC)g\/fE6fTWCd8H?E5D4T#AF?7=H-4_:JQ5SHXa.7fYMBTUIMVE6:+QF1Z?
F,+ZQW+U5UEEfUILVU?;GCGOKR(X#?.Ee?70NB3Q3C)3X98P1GR6IU:+@c<DdC[_
1]9A(2]Cg?.^<?WP92c5U(ePJQ)58@LeP3Y?+;F46JIg9@6BK2b3(RbR?S6V;>@M
T)[2=+Q=gAVAX=V[\AaV<J&@g3GBH[0;5TR?393f9X+eN8aT]:,VYb+f@P_JR3:M
;;b,f04Y(f/R,4@7AIDX-:<BN8SKbTZ;KP=\gg:EPZX8[0A6.1D#P,I?@K:5@d_8
)8;Q2[Lf7\HHeBKGeW95_[J@N65[WJY8YF)a&;Jc#<@X&3R7\gb989P:(V?I;Me&
QQ0HH2G\_ZW[@-5S8JL.0ULgY:1a[YbT.4+\&)064CU=KgVZ9/TL3AFX14L+/I?4
f39CT]V9^TJYSWM74A7R[D0G4,6X:c<L9MZ+VHKf8E91,D@;2(3PDX54#>W/P[^S
HK.g;@[U.cGMML?AOeC/0F)@CMO,UJ6c#N5HJ#8R8VO:(ARd4D(g3-5BFLE4T8e<
90XK\F+WYb1(9<dD[\HZ/G43I]G6eC;L+BSMV?3,#Ee0aeQZ@^gK<CF2>1VU=PcB
?g3+c)3YSXLJ=XgMFM[&?Dd^O>55@e?^B,b&[Sd<8-7Z35B29L\H+Q/,e/S>[K[/
XH[T;[QBO>7WPgG).<)WMRJ>_CT,(I^4@0@&NF\?+&d_a\F^ER8HK?@[U>Z=bP2P
GH0b++T8?g_Tc^>\@V93a#O;2IGMFY,TNSe]QCZC:DH+\b0N@4CB9WT8]0f-12?L
aBO@J/a_T#:GTJ^=DgQ3Cgd38(f<T&_NOWFb##AA;VG/-D8(_@/^2cKG-48MfJ_J
,>3f265Da(0I:FW4(L/SU_P.d0MDYS<eZ9=)fYDSACa]fbU:4LT-DNTM?CC35F3N
fYB/62I9D4\F61\G^2TZgD7c.dS[8L2#YYV+:B/Z)L0JfO@]Q.31@0U9g&#6G+U(
GC2\XINL^P^08[ecR,e1&;MFEB5U9fYFI4&JXO^ZJRYL[+S>VTYJ.dV7H=e51TZ)
<E:5G=@6-];PF#I?TcL0Fd3d@GgCfgN[LU>]eOS?Jg::<fcHIXDXg=#]W394G[]0
G4(+5f<B3]g+0fTHA.W5H<Z8Lb5OXaZ[MD8NIR;K3Ae(0#NScTYIN_De=NfBPN87
NMDbg#b#[HIAEgJd5>;[Q>5;>VKE1,e6CM1XX>GdCb^e3V&bW.+Y,S_)Hb&,T\XG
P5T)PHL?@7-3?IegZ22S\&]QO+@0SBW7NR5D3J:]2,XFRWZ/JDHYI_=J53R2J(Uc
^N\7?1eRS0JfXg+Fb,,9KY,JeUN,<4]+EUTa/;[\5gHaPZ.dOZQPJ)e[QcSQQLR2
NQHTQb+6La^@eJP1XS&G@Dg5B2)+BUf]e/0NIV9<6C2WGfTZFc_-6H_196LT1g.C
^8NY,B9LZ5a1)@ADVPV6+.L,0J_)fN;ZET]aLEM@&IeL5)DIAZUF>T.Zc7]ZbQS=
>BW:;5-:UOfKR11KD8aV@VXa7E<e06VdTX\NEL[e.c>[(d5aa/&f]-g_1A:O2JQE
X)Q1I/G_FVaB/9Sg?,+@1.NQ/BLE?5geD9cA9-;Q#/+7G?/If.:VcE._)C][BZ4.
Id#)D+M&G4,QC&LU[=_UVb12X26Y:==5X?C/:f((77#7_-13XQK:Z(7ETX:Jb#T;
A>BC8^N>4G3-_)8N#Z2NGJ[D4N)8^\TX93VAX@@Kc/YC<+Z,-e_,bGbG27\YD7gK
Fc+(a39BN?fK?&UR(C;\B(c^=L(@D+2/X=J2-\&VJA(,+c.gg.N5Ge33MH.F/C,,
J9PbL+=D#](#^B^Y/1/0E3:N+acdP&J=a7S8JOb&9BPQ_4BIOX[Va^R3-\[U;c(+
N(3/U/,bNgJ^L&O]15Y1c-32I\&BEAc<;\8<4_;-WXZ&+CfgI35UD<2N<I9&Y2-1
WL#]_2gJEZ\g9)B3I0^,I#<:2+EGRWf@9e/(Y/P53@29GYR[:>g[+8UgG=6bZZSS
PT+GIDgJLXW#,&E8SUGf17W;e7+/9T62e5C[+Dg5UU?&dU5ceHL0NgfQ;)I^M=gR
+:(WARB#9e2g@&(U,;@@:@=bbaeE7M,DLcF:<U?d0U_PW8(5J7S8a&&[?FQTOMKX
^b2DRdgMAW2d7>AV6>GA.::K?R)c/7<0QK=)Ob<C?>#F^XbH(E<]3.CDH9J(8b_Z
I)#]Lba6_)SA+S5#PBLT79g=7-2@L_<B:e[LW7M)JMJY((KfXFASVT\cQE[B#TDG
HEYc)^ReWIRVDA8XB,RX5EJbGT4:L?g,Y8Hf7^NG#KObdK]8D0OFa#=V\,&QE7DM
NX?U+A;a(.\B+EX-d-WJ(IeYK(5Pcb]XN0XOP+/Y\K3Y.)EdT7]f=/HBZC&-\=4V
>f5M5Cc3>4NXHKE.R[5)FWA8T7#bR:H:I96KDAc3.Cd#bM+#P0/_^F/X?S6;V=RK
3^N?S#T3P83SY5_#0LbEB-e@Jg,1d==</LK=H-a@;VF,TgA1G<+,@MQ)B)IIP6-c
UMO?BU^WeCK?GA3&.[>G\L0_gW6:L53B,,WL:J@:(I,\[YaE42RI9WLg062eI[-M
JTYT7O:\3#J0BJZO@gUB&HHRRA5@7ecIX42T<)dM^<,Z6&#9YB4>\.e+a0ET[=?W
]g4QBd_LU<T<K90a?NPI^;P1J,aBgeMUCS9:#CIEG;TQ^5<ZQNR.E6D3c=Y)[[a<
@Pf-L4#U0MEDSeW^^]K]CX8;\,.@[H^8P5[M6(H3/90:F>+YFHYR,b]YFNON>ZX,
]-HTSVYY3^=AcGQ/+@#Z?7cVW&Se_74KBe+),CEEX]I#g(bf:DgQD>YLR6SW=1R.
ZZV;7H:Y?OWBSTKf5D;T+FR5b^5b-P)\<S\6IR9^LX.G(^fMJ@6HUeX@Y4<JZ1SS
CPK&#GF(3Tc=,71.)[5^\cX\#?:\99.2dV:bAU#b]18:HEFc[D3Sg39S:NSc7/Ce
0YZ,P+(J^0TMV.P1<Q56;f\@CCW:VF>KC[9=CMN7[RL]=D]+A8QWR#ZIS]M^ADbd
IbHaER?WTYRaJK>L3d>YW=SC9AF6C^XO=L6Y]&YF&W_H6QK--CbVBBN8;S?7a3]f
W/NdJ__M,=5Q@8CK;6EXY;V@B9G9@3QQ0d?fe1S816]1_B@WW:Z:JA?&(-2DD@^B
_]\7X0Y,<4ABPO+?fN4<>;I>.L+^#.QL.11L,\XB,N>;GQfVK@JP\WOI<<K8OL\c
fHM5Ae.,e@3ML(R3WH@C7@#fg-00^cA2VTU45TB3\BIBE+CR6RQY_eNcAX1T,2-_
^<8=&A+f+[:H3UQW(c#AC]-ASUL0#McZ#OAA&5&aAZ=g.Yd/XDe\^7#BNT[9cLM^
e@eTcZUAFIa1X=JYY(_X<^_J6_P\#JPRgg,Z^Oa.;7+BfOO_?Y.:0ebT<GBU@4].
K?DQg-Z33[4SF,T=\2XVLcFI+:]WB,)g?2;L_ZQX&<\5R)FM-(K9L6KO]dB4)Y^6
C62:9XE<UAALR/CC5)<L2E?J/+9_g+1^bZLQ(]TFQL.eL^La(C#C)XHVQ7e^>gL)
H7P/6H/DRSB:RU/,_RPS\WCYEDQP]dF.S_.[ZZ.HCbZZS=51T43_R#e2Y40^+M9<
I+2^;#:/0f1L,.:-]V@f<.S@.gLCLF_#_Y1)C<cFCC#GH#NPa[c-=gIWHGUb0W]#
ZZ:TR3NQ5O-f=ef>NJ<+,15\#YgIFaF&TR;\a)ZV+DKZ&16PeR3.:JV:3e7c?32^
E0XX[:T.T:(+#T1\#?:I5:F_@3\4D5X&1DN_O7)@;P>G//T_eS-A.H0:K4VYZcIT
:#Q4C1VBKc@,077LM0BY)UW;U#<8-gaAIIRRZ-+L9:+698>.b5\8(3LIC@UgP_)T
bIKE:B5Q&S)CT<g_VZ?CgCJ9J2IcEJT3V6]X7VNP@@@K7BH_.[IJVIRc]Y[J.XN?
4K2)9-A532M;a<0UOGO(1Z=bCI6Yb771^NNI,g^607UNWX>9]40&Nc>NCYD-A8Q/
ZZ[U3R:<ZVECZY_<7V/QcSQT4NR&03c]JGH]ITd7AD@bPG^N,Y/5P3XJZL3B9+]H
)2Q,[+U@J\WIBU-GPU4#<L3NWB2QM@e2?M#a]FF?<Za.41M.IPU9)N_814gXLTTE
cTaSVLI@X.7HgY,EWI=PE5QdT)+Oa]d7ea4XQ.Y[RLg;)PdePXJ_cRFSN?J2e6D7
?PWRS2Sc:28FdaBTPQ3WdCU[N[[\ZI-]K@^Y-OQNJAH0_T7)W_#Pa<DDQ=[5C447
B&XBOFUK;PQ.>OgN,_R/XG7(NG#fZ3J)c33DC,3<>8K@8CQ&:@T9M@6FB7YQF\X#
\<80U4:6#M=&_(E_^Yf?LXQX)-.3)[g-:DL\QRBOV>D0UQ;eSOAKBeF9:DX;a#6^
cb@86]_CXEPB9IgdBIR=+=UMLUc9V:V>(0AF7af^F4GJ+BA>#5S@65O.2Z/Z#>_E
=YY=:+58/B:cZKR]-6>IU;>KEgWE6O;?5Q^@g2#[G309^XTWGRd@[L2g-9IM2&X)
/^74bF9[C]Z>Bb=/?U:+d(_Ka3D8.X&&N\0AHeJWPg_?>(3DM<1gC()&H>K))S1.
Y,H+c1\Z5>5I,XX#&UN9R]-R=R)AJ26V-YA42;>JAP9LJS55=G?GG+5;acV0#=#@
,dg^Z1^(8;5K3>#)<>g]Ee\EdSZN1.IK6Sd3>-TQY(.eW,FaC[VX97WaN)II=P,K
1c&&A8/A(ZfF<\@/^DAY4>7/SOHbVZ+=,BP&Q8<NIXZ:]_1#&F=&Z-20NLcQ6]PF
6Bed6#&MLC5-.W688D:@N:WF##S2b?5CgN@gBb^4]GY]a0ecQD/0B+=]TGgYQBe@
5&;>CE6UF_<-J9<QCVE6(H\3b_V/H.&/U7NSEEe&:A1,_C9XCHG<AP:GJfVcXI57
JBZ>+ZZ.[#KSa>I(B26D)#15T&e=^a[+8HDRcT@Z6><;<B1AcV15<(VL(^=AL+;&
.,^1N<M=9)2I[K+LE_I&ZTeBW1;67N91:d#12a<R+CfQQZ35V55P(eb)fN2)U&SA
\/+E.L<WFX1CO70B<NBGUL#::C6[bO[5V6dWH,Ef1[Pd(87V,S1T:>;Vb+VT5Y@D
#b2WfETgG8Cd0/eZR6f0#]=?QDMbMT5b(Vd.,2Ae2U_+@1Z(?/fDMZEAeM8IN0Ge
:a7G6K0P&/>5JA39.g0^MaD-gE#gITBY5FLg6ZK:#[0FX8cIA<7MS\#GEW.@3eAP
dO[6D/g@ODY.T,AF,_.;dc:54MRE(MW@P2]]Q:\J?d4:I9gC>2)<L(T83J^X,1#6
CE\4G_@ZbPJN=7VQ=N_E:c[Mg9/905Ud_f,N]d7[e;@NE7&SCCc0;T?/UB2LA:QS
I#8]:ED:Kb]28Eb3f[W]U^M]QeF:H#BIIc+[;7;e[#&S25+e4)UQO?<F/T@Y^Uc>
@>G.6N&d.a2U<Bg\,0]K;Z#7HH)/CbADa9Ef:d)E]1C<PS.B)e#L@B(2Q3XCc#>G
2OYJ13CE-2V8c1=6B-eF/=DI5?N]9[].;(_#((>c8]+8?5;d/\<3_#PP=,CBCOW[
BQa73OEGH]bfIS?F#AJC9A4d-6TfZRB]ME4D[55eKIS._90/:5[/X0HU_KQJg=.3
?W[5J>gE+U9aZ@/c#03D]HN7deGBGJfg4cZI10B@Qe@?-G)FN6O<;VU?b[da9E:8
AfdLRZP^PKM>Ie1[EP[,_W--EE(2?,(?fL-aB82cO?1B]8,GH-V^Z:Q\3H@LXGYF
8-Y4_2F87/?bT-D8[>5Qf7JHL:9Z=HgIc)#^851XSB&(99QLDFPEEeA+VfUTS&Md
d-&T_UP=#5d_N7O,2(])Ee;9aHZ@7L2,)3_BYK9IQMPfTW\8KaRe8Q[0]YED?M.8
bSb;?f;OKa5NE&T#WL9MHG]C^f6LP=77LeYLORQ15:0#./(ZI7GKeT-E\aSaV4a]
Xe5TFMZ4]:GAfO:68DdA/D=ZRa\.49=7&[)<;NWAC_cb(&IT#RJT5E6NdFNRFT\?
DNKWPQb^7#KO>f-Z@?-9TCB9AJYdCE2Y2[ceS274#82ca&QRL>HYW]OFCWS;&Q]O
<<M\WgK<ZNJKC&5#F]9IBGeG;..2;E2#D6UYS/T:f\Md)8\=IKFRC-REC^@AGOH@
V5RCe7UY)K9RVJD:(4M:L8+^dC12TO29@ND?>#TRac,=+?VQLN3&O&XP[FK47=21
)]KRUI^N_92+>OW_G^S-eHGCN+f3XJ<U-.GgL6ce5OAV8d,7LNJFb^<N(D:6(DKY
P5H]IA#.96X6#&4TLdV?aVdAE1A([4_1&+X\3V_MI(<3OY^a#0)S2.98A0K-(GN-
ZNe]D5Q#WTaS:2DB]b9RCJ)-VW0dQV&>F/.\9NQFKC>EG/(.@aI]LD2<1HX+(@<8
0)-a=WQPDTbgU>_9d.8fEb8LHE:BM50J)T(^T;HVO99VP^N8cR5dEM9@81#5d+U4
W]SF7X5Aa;VUQY-D:N)&+;^0AZW622Dg.4N>SDD/]f6+OXX<-?(3_6-H^ae<W=cE
@Rf>6/5CNeTO3P:@gfDEPb)>65B><^5O70MAf+.?LSb_EL2B+@&I0SEC[^>b==D+
Z=TO@&EdK2gBL#TAB+e9J1#\aEN_\F,3g]d#N7Z;ECaC/^P8c5)_Q8W&R46gaPY,
^]0L[./,7IaWDW3a4Yg7I)84>8-IIFWT7LQZ3-Xa=Rc7CTBN[<NHf820WfD@_MRf
:^Kd/6NRG/-<,[<8S#/6)Ye5OL:.Kd[EN1=M/TJ3YJBg1]0e6V)>SNNa_@gI-_,a
N21cWOADK-e6##6BT4^X+8BXdXQFI]QAPUM5[)V4f+fB:SBGJJ3BOb07/@Mb4W7b
0J6IfASed/297-Z(O2]#Q>UI)DUNU<N5MA#^O_3de@B@QITH[4=W4dRdNZ^W.8Ia
d&8?gC0AQDe&8#fE:6I3JI4?&AffbX;eX_C?P]cH=#4:K9-<7/]33<2JY@+V3a@c
6L:?M]7?U5+20M_#TZ(B]8]fHGV=;#YgQ9VJQ41G[PcO7eDGA1@>-/>f\;PQY]5S
F4/VDf:HcYL^L(-KT^V&P]QTX)<&Tg12D.9-_1ZOPK<ZYYRKW2+,f\J+@f#g6V5D
KR^Q<;LVD8^U?;)EL__0_SH=XWZ[U1QF3.E>HFPKZP15<TWZ,1AX384_4VGL_\&M
ZW(LRe1PLRY@ZF1[Dc7\@eJ:FJ)Y[GHA?WbGI=([13Td>+:32;AMdE)[]H]XD&OJ
[b(ME6d1T+TNK/?>.VA^1WDY2]DBB(N9e;eN4GQ0b#:g[e)<NVA+FRFa1^4Y-dA&
a&:7bNB/@FQEQYa_&1[WFSY2K4TPcg<Z9RM+M#:a:/?B+.#fWHL.39\]Y9?C>N.g
VHWb,9002]?A-.&(E#WB)-.gLY0b]FJGNIT38QeA(25:fLaMOUIE&f:3H5Fc?2_.
#7&;H];-)YNe/-,J]dS6A7P[[(U[Af^)C:MRP&6eAC1.G382\=\30FLOTBV=bYQ5
VZZ_Jb?MA[EWd6a1QO<PYTY@8N+KA6,CN18,2d3cXVI3gJ[8=0-D,K6E941SEX7#
A[),Q?5(,CVHD080+J48]I8#,\XfDZ258c(-VXH&[QfH(.CHD39S-Nf\Q8LBfG[M
T<#LeeE#4]UOE^Zbec4#ONW&\+0=.gf3:\K1E_SdUI3L^(F0&_K;I:dVBN.;N^Hb
ba\).QO<&:?3]>NK9C-EUG+T=C]Zc=fWHLUPX)GRM4f#><S)NLJ24&c,YceZ=W)^
aO2;L0].XSBR?VL[cN04R=5K#9@RG\Q(C+L8(dDFYNP_)]]2=b+J,b-T^0+dN7OF
>F@bb5QS/])SR<Z2EEAP#\CBB;ZG.BQHcKLF3AAAOb?AB9>BE@7Y?R8a3;RfU6FZ
QZeG(6U,9=L&SI2cYJ(&X@dRF3R,9M+Y>&R2HPA&/Pf]a#&5;74_BH->K3C&JURc
-Gd0?J-Qf#PA8UV,_=abfH#6Pg^QP(GVTP)a##ZVF5[5g.fL5#M9ZU_bVH<V,eg:
M2R3->DG6Rb&HN1;36@6PR#KMH+E\@ROeGKR8UA/d;TaZ1K(Ig>,F-=OS@M<=STY
56TMU@2+LLdY=/=DE_@W3V/LPK7.7;C>=A;U:[NYD;TWJTMG]Y0M01>:ZYbXN?We
GDbd:4_HQL>P\S4.:4YDeNUC0L.H;[>Tf#-FQcA5#+f(bfcI.M<R6J/):c<d:>Of
,D\8ff/8L#dCL<)(]K(83.3LV1FW>a=OV)[C+eII6@^Hd1RgTP97bN#5B\HX)JX/
E79Q[=E+A0TBaMH86eVXg2,2edBZI[HBaK,SfZNRI@7;CZ8-5Ua#BK0;IU@B:6S]
5D0:g@1Ua7e^G5]&QI:E@B24FDUV\T?TWJZI7Hd#YM0)A8C)#_KB>HaK2fOEd1M+
-=8HbQ.fKEbf],9J_L,H3gTFN&=\8]G.;bQ>(Hg92[#WgZKc=8SPW:_U81A33>(6
=/X29@UcOUg)3[956gR,(K/1=HHZM93DPO>1?0KZ:B&I(dLJ#)^ag9DTZ.[M8(:b
Rb4X^2ANO<).gDgYb7Jbg52B#IW+DcEJc?YX@bI:Af0D;QII71:UZS31W<)SHBX4
(?(G-a_B([GR[d^Od<,/f&eB)UJ#f@)S,_\^]2Y556,7OaZ:f8]60?gQ?G8d^;WH
EM^56/QDD3/VM@5OG(>@b&dO5G-3\4(LV5aI8QAPJ_T8@--0J9>-;^4Ka7^55ZX^
@06X:6/8-/SVT]]99EW:)#(Pb4gCJGV449ALe.3O&3,JH1D4B[3@E9K[:NEMADdd
9E-0SJV6C#@3g;UaR;.;>H(L@1T.D3N>LKI6P+<Cb6XPLZ#UW&OZ-[\[gcFFgNLI
-aebgV94U>^BJT.[C?A<E6JF3IS0b:JOP,FAUAB^FT8#)F/<+HaTS/W&^#L&-Q]N
Yb3Ic:R[dF#3K[0V@#A\e9YLd6F=Nb+>7(R:O3/_V-X\;9R85.3c@K[M+36QC0<a
-fR(Gc>(?.?@)M:bX]a[R7(]6\H=5L#ba/;;Z<4+g\P-HSX.&N9TbbL22L:.=SA:
ed@-[WG2gHV2+YPCWPI-PNF)#Rf1@@>M.06&M>D^2Jb^]333(:ZPZDfYLCNce\<#
334gAOW=f+LVXS3DZ42>VC62Ce:,X]U>V?CfSEOU?CHPKbZ?)KbVW.U>_T.F#TdA
\N>NTceMe7CT:58:-/d4gV/AFTKeaQ>7>WfVWEMM9[UG_R#W=L7\a4dK19G8YR1c
ee.2^P_?[^YLTHJ@&R1WF1bcabfM=Z3L-)L/:,Z4SF.[fdVMZf/QD03&W0K_1HEP
I;DM=b+]HY?J]cU]FFB>K\,<K6THf=Qf-gIaD:21XVG]WNC>>?gG6INP@FPQFS@/
:=b=KFRQ4X/=H.9HIcPZeG2Oe;424DHZ3WZP3dLTC=JI\T4)XOaMFIVJeVe]b^,D
8g^7Y];;D=:J(Y[[=>0-0]/M=d[[JA2#]?e;,YTQ=-^VH27ea-+E#GHa6f6PZBZ[
7[eU,]F:B^9><8RMJJHdB1.>,,#:J9H+)HI]X;=W,gUSV-P-)R0ZX=Y_Y=,)YW31
3/M7KV>_&aZYYUF5?9,\_PDOH8?D\3YL]c:K8;G/>QN<D7[0a&Z7W&,Z)U\Ng<@@
_4URF6c+GAW2>.O\LE[-aFA1<:QPZIb&bYP:Z4<AYU&/Og]D2?[#O-.&;9R@?T]Y
&FJRRb;LYa@K&UX_+W&SeQVA^cO<UW;E2A:L2g(C9JQ-Q@0;7>\)Q?-&8YR=UCbA
:eG\\5_#]:>G)JRI#P/GW2IMFe@)?CAR?X,(ege,Mb_f3-L)^N+fC_QX#g#5F3S;
A3HCd619fgWFX72F^9RP.OIVTNbDM,GZ..cDZ7_Hg_Ib6PK<eFT2^[O=Y&N^UfLf
Z7JebG=F=?f\G^]^)b[CVM&cY84KF&7dOSD47\ISQK1TY#NR/4]KIZ:=e&9(92@0
GFb.^H5U:e382U4+g):V@^UEb(eG-1:GP0^Q7MR2<KeI:OR225?,B?d3_.S,fc?8
\F(fa_,NLb/9d/+N\X;YEfEgUI6Ie;Q:D^_<<2DWafUc&=c\[CcR@+7a&CWQg4?J
.^9^)G5e3(2H(E1P#+PJD-;PaCGKCKB]X?AM,[eDCJ:6ZT9Ycc?E+_,5c=f+;g3=
HeJ2g-+ef62I7a1JG6JN44I)2Pc>.5_15gH5RT4OO(X-@WbWN>3XQ;[a0G8/.aID
8JBL5+EE#g);3ac-#UM1Zde@+aO#L_WZ(&Wd\(#,L/EN?UQ10QFNKaFLE).1U(\M
Y#\gET22,94H5(cB6R>NZ#AT/7QOacbD[Z7ZEZ\gD@JMU]+T68/-K)c77,e@aOOe
JdR+)a&6UWGNYBD>Qc&X2B+8:IUNF\&+bVS:f6:,.e=;T?OgU/^=BH07Ba>CN(>3
)O7+^;2BC#,8cF1MLUQYM71?M^IM/AQZJQ2JC(c3U_A-6,ZQ6Z_0X&ZU#YW[4GYY
;QIU=\B-T\0?-HEd9YYgSe9BDLG5TCYO0cA?=A>04IMZ2:_I.(ZML5:XBg@P-XR@
=SF876.9JI+2#?LGOD@0<ab&c+Z[^<P<:BR)WX.a-;f6-Y:0.T4I#-8?^68W/_HE
NIb<Z^O<;)98CgK11&@a2[6P=+N1fNd<^C_84H_=]Q9JcQBW7@(+=e<>Z+B+#H32
[@T>dAQ_UTPcNL&)/bG#Y=&:e3Na;EO)-02K.R\cEQ3bN[];(:fEP56U.XL#A3YU
4&+1=-bD;CcbRO+KMKM,(SFM0NdNGV-&aFW,5[5f)_[XIX/72,P;B+[1I5^X#/T-
dN[b@fA_dOQ3H)SdVMT4H=0g7>9e^_E0KTBRSJ/gJdfQPeM-4L-bWD=C-^I6cKQ/
:]9Ea]eH&Z6O3+aM<FG5,C\_-;W3](ULcYG1D]RGV<-MPFTA)6N3A\5EV#1NNL7c
XPA;V@R0V;_W-SaT/;.PK4U>V]A(?eGLRa[dLCZ-9T>bL(]<FU41]57<HN.0PVLW
M((CSXcY-^85g,_C@1ZU8?\=OS?]]/33,[,K1W7;;fS^_We5/-ZcPAU9<>UbS=S>
EKb>?\aZ\9Ucb#X3UC1/,UWSM[JX,-W3bMK]g[RJO/e_5d<SE4ULJTW>+U\8GCC#
C2-\0.LMDIPWADe3L_P(_&Y<+_\7;f_M5##+W;S^N<fGURJRD<WT?g00JVWbXUG+
+W39#R]I^U+H./RV7.e,I(1L)>G+V]I@H0?a-H0EZU]VcCT9CZgJ&JNJ1GeSMJf8
#]V/>aE_&#.UH8Q@NLT1C):CeY4WN?9\&DaQB;W<C+<^6BF:Ybc=350M&[W^6fFC
F4X#[/@KO#M+^:6[OR#Y.&\54Ff_4NaSdb8VDXGE7F)e<QN)G:F@dXK\LAINA2J:
-c]f8&geB]<,-A>?#D+PCH\MW,D8P5Q3IX(P5#MH@Ge7TXLY39Ibc9UYCWK(N7([
2V.EB&UeGU;F+HIH9.->375VWScTQ\3NSSXU.1eeT<;KPJf@4UAGP:Q]64YV/PfU
ZQ@f^:Z1#XF5JL?fe_(X<-BB95FGO1&:_[::@ER.\gW/GV#G01PZBb<H2KP3)AX#
@9fKW7@7H2UN./0dJLQ7U#L&gJ2D0H?GgS#><0;f\e(?XaR),>U^3KQVPXS?&E>T
;I;&/&<0)02^(.TKT\YI(W38IIH/>;_;?g8f37b2.]L=fD.LPMTVB6_0NGJg8BC6
e-b@[PbH,JZ>]<R5e.ECU?X;IXM5(V[:g^RJ)]XabT-L#cCJ>[RdCc<X7MUU+EZ@
WK0@bVI#<)d02fA3:>VRPF=a-3SdgOWSR>12?MF5^3f)94/G6V@<Z=48f:8PMEVL
]T;GO<(B(4?N/;-ZR&_X@C\Z9S5c(c_INC_YaacX)]M=I)G/&V)TB78D&@:b,HH#
[RS?89d1Je8cP,/#-7,6EVVgXJ@[bd?@3eL,ZEAd5PWO9/_I?MDAQV+]J9L(34\_
eYaIfRUITKQ<.612I)(8(^KC^W2O7(VBd:ZH(=FB#0VbA/23@Ac.Q_0E[XQXFXE)
Yc-[7K;<VNBFeW.FeJ/YHA3@>1K>;5PK7+4dd->7B9-.-eQQ>N@,(IUSI=YI2HG5
\EeVJGP0T>(KLK_g5OARKO>L<>VYS#-LQ\bf,1N3^7e/cP-(2HadeU[NJ\(bTa(^
Dfc);TNKg7T4:8,M(&.](7B]PTMQ^Sc]>T.\XE48+7I4L2/<NWC(g/Sg5)]0G&.E
VBU-CXNOVUZC2&[S5Y:2.Sa^7#5?WN6e+d/YPU7a,KW42WZ9;PbU&Z#45-)9HR2K
;AD8@J8/.)=aI;;JW9YdAa0Y+;P)_@UCS&>P[Le5f<f)+L;b-f?&g9[@VT,5feN1
D0[-U&.VK(<5810-X+^B@LVEdf]#2SA&\<S@[^J#^V55P(P9D:aHL#NG-JY+Y(b[
LKBZ5&OCUW4(\=+?QNSCP9a+e=END>[L5^@0V_DO^=R+_3+H0^,aQ_B=YR-HFMMe
[B[<15YS0c)E.LgRV8aGK[6FGeAD,H7FYV<H2PI\7J+B^V>F\>_A\\GUaKf>G0+I
>R)HXV9;38S7B/EZD&2L:TOXcQY(LV-U4W(d>P,:9^eX&L91Q]D<DX/P6G;cg07G
Q,C5/.(AP^?Y>K>c7,#cEe)I5;#DSOcTA?<X94_I)BdQc-RN&>,F7U,9A8af=^2I
6\af8=<8[)BWRT9#d9gI,Z>@9BW^P<?_HXbac<?G](39:D-A;AE+_PdBb?I8M=13
;^R+_KUF26?FDEW/]C=@C?\)SVMQ<D^+gd0#QY_b,Gc-d,&K#;#5@-EM]@Tb](6V
D4_d-c;O4J/DWH24BQ&1E9TK:b4YX2<\b81.?\TK<\@Kb_LCZT28U]GP<+IZWW][
&F&FbL/H(1NaWKU)VK.Q]Y.2N&WeTF-eM6F#_;-D7:/=Gcdc[aSe1Z@#0]e51U>#
669Z^L9MVcdc(6eTA)9Y\;<INN&+(U7AG1FGbPe_fQ#.>/_ZLYJ<ZD3P60.^S]dN
FBRZ42V)RY]K+I^AE43O89CQ_=9XVE,4dQ7UC;CZP9aYP,>G)_\dd&T,Pb]ZgW@J
-8+TO?U6O?a&)HJcVOCBTC-=.U2G3<V?9F^)f]],6cKY1EC\O^[SG@3-C\W/K(&,
+T:P^aKVA_K_E=EX5cN_T<G(CN4WgVVe?gKS<5F/X<)6I16TW3GQ+V,FA6T>^&aR
\]+P\:6PU8=C71#B]X&MKV196Q0:#Rf1]dbgN-[Q?_SO;(?QUQ?>40XLJ(:TFKSH
g8=G[_6<K=TE][f_&5\&PUbO60D7]0fdA_BS-=Y_S&9@HEbHWGM(F-7c&.CFK__T
>SSV.2C>EV>8dc<#&>YVDe(BNb5ZD+3,1689+D9NJB=]3&2LVKI,2^I//_YfJ2cZ
S0RgV1aU[LIe2E0GQ.(X;>:a(>RUB95cOE:<edL4Q\QgJ7&,5d@:P+YKBaORN@aX
DJFVA2:ODbDeFT<fH@HN<YN:a[)&a>dZYUH7)C,TZ(57T_0U]J=77DGK7gVfKL]d
\=B;H=9F#/g^9;44fGTLED?#T8W]G6PLU^UVWXE:9L7[M0KE,=T&/T?>Z+1,C>Wd
@-48]-_[8#IMP,<HcX5E.VAaZS0U3Y1O).B4G70aAHJ;?5F7J):S-c9/6[O_ZB:e
cLLH<eXMD+HJV[_gNed.O>J3:b-:L.-AN?4U-W4PNZZ@:;_0V\;XIGB^b;]:/76+
NDfG?T&dNHMT9F[f&/5,[F@?Z-AOUV7fK;[Ib4PXQ#>IV,1IO]5:a]eGKO@,I&\=
RD\cXFe)>277?+5:^^JT_KH(JC>M:7EB+WA2/.U&;MAZTg4Q\GJI18@/8[)A[Q#D
HWQR8e6gVb3P>#GIbY)Cd_<:]eNDB_-aMV4@08>(QE#-/_VL,c3EPI<fc+A_fZR@
-P#Kf_@H?g+<M&-GFeM#KDIQeLYK?<UV8,8d)F2X2#I0c8FOO-4P.T@U=5FY4J2e
R-DUV(9(U2/[5@dg1ES,XG5OYb>A?94C_Q+?OMYYaca/HXKMe(GeG<CW0/Y)C#e;
QPDN/2-8Mf@#aXU>QJ6J>XOJNG1CdKB(fX3f?S+#f0g/Jed1N+>-Vg.45QT#>0QZ
@R42/HV8c4.PXb^J=M.;FU2EFZGd>&VOZeI&#DOEe+DL>7^PV98O=_<QBJEM=JE;
AY4aFb2M)@PaKD.QY@-aOdKBP_+FB3K,<SA2Z^:-X+fNg..FO<Q-+Tf&,<.QS(A_
H;6NML3(cYc/,;_TI=I0UOeI34LT)^YCX<5XKVXG<^>KG_MGZfL=g[J0C_XeH<eQ
&eAB8(T3T+U4H:dd;YIRT0]c3FR563_3O\Q#2R0,5JB.KR62Y#0g,>/G=@=L2T=f
[ea1_BcV#H;fH&L32eWWf07+WJ_LLUO7g<,TM#-\[5(V1#L5V3F:#7ZBGO@I4ZZ7
#B(UXU?ZWg6E)a?5ZAPV2C<BC160UZdbBDV:ROKM_]\WQI?3#M1W.X)gL4G;5G8)
#G]4=D8QI2E2EX1UegB1OTN2XH&_3S[JU8.S\b8RVCeB2RU4_.=+M^I-N2((A-DH
e/,;L_d=[5G9cI6JFQI3)fAaCU_<;>d5&8U@X8O=\e;9#/=5-S=T,g.a[I.eaLO&
_&_]7EL7X=1W&LC#SF-)V=CB+f_NPWKO-<9QG7Ze;RbE.82f<g#_XQ9CXB,d@8G1
<QLX@>JZ&2gJ]#9.B6e15+D=7]SDcSX:^\;YO8\VC^UH/a#7J&E3aB&dQEL?WUBT
03Q.#F3EO/d)[5.+<<3&^_\VJQ-,#5(dL+4/ERMI;^U@[=1>T>OOYX(_S(IEeI5B
A(9^8dS;DL)]5LI\@90P[,:Q9E3HfD:c73g)05(7_#R94?>5Sb,BIbI[P94cO2?.
H.2gcXLRUES])XCUY59gbDRKDfI1HA^cZ3V2J0B@>Q0,.JFfe7)KW.H=WfV.BC]#
J^O^4=+b7:R)cN#0Q@4-g]b;MT2#],<M06-R(\IZ3PfRbWMQ(ERe6E_EEP\2;O6G
@5?VRZf.6?gJ?DRWIDTQXOQ:KfOXY=3U8BU6[,3dc&T_eKBOG)#68W/T?\JPI1ST
4[EO4/,<M7AOI(@=C>)2-(E,N.BEQe05?aX=B(fAH(_X>Ca8bW.5;995Nb]+X31+
TR-fF6H/2TN-b;;X/d3X2UKXGW\SYCS^(Xd=fNK1BJ=TF_?Q9Ng/bAgf^UN#0U0H
<:^EAPA-F&LD>Q:FYZ,U[NI^1O4(]B,cb-X^=e1>12@6e?cF]41,K-/AT+,(/0Q;
LN4@.;O&\<QMR>NdADB3CZ[RB3M4?b+5CZU2cZSDLNg6MIE=fX:J[F.M/^U,d?J:
Ff)@.<ec:=[cSU,;@>[8WG?OKS8Kd]Q^V@<IL0+I<3(1=.egJ>U+Z2X-JcR_(:^1
(DN#6?ZeCF2O;\WYWg&M&:SC_@T]D?_)Y9N1_W8PX+2#J5bKCYW_&+UV=,a0W)<1
P(KV2IJAL[-XDHJQ/EB^3_d99He-=O23Md,I)^g9Jb.-X+J=CaOYJdGe#Y]NG3]@
JP5@7bR]@&UAF=>.<d-I1df#IGd4&]eUb26K=D)685_>g3D^(Jc46J)fV2b\74]+
d@Q>\JTLN+OdZ4H[IH,RP1M<08Y.8gS8X^S6A.G^W2R&0^YD-FC16J2JAPJfNgg8
_:YF,^\a@/0)^OW0UYVAd;;H.536/HY:];f:USSE8O@&&([M&X/]bOAE1WN)6)X0
Ff98]E4Cd;+[/0H;FJfT&V[RJ7_=6NZLY+/B<:59KfEZR&Ee7O@-8f+GZ4D,aPME
fZX\c?L_@EJPTC^\#8b5TDEFFSO^7:B7c#Y4=;PV(HZ=2D-Rg;UZF]\H^aS](?9U
07=YaAV;N&MU\]+NDKI[6>1Db-a.9[)[P_84?=G-++0_I#_JK,E7I;3ZIP[0,<D:
PQaXffZPN/e1U_W8/]/KB0fMgH,0]/=+C;:/Ga65\O<_U51:PT4(.2>d<E,_(Qa^
L=;L=+0._d0_I0.EH1^=\,Y?2K/S&T_#Z<(9]CSMWDZKM5]WE&GEH:_Wb>>O#(b#
M]Y:URfOX2L@?20<NWc1&W6(&^@MT_1_Gf<T._d.5744T#OU-+Ue2a.9:)+342G5
+HD]f=JXLAWSK+W4Y6bDKQbFRA+D#.X[e)//B],/A]O:G8DB@Q;:#0DKc/JTH)=;
(Z^([N.61A,,3YC,GQR/AL?6Ref7Z@-9F\L(a),PJ<V)P5@+F1B_,H&cCRDRW:2P
P[2aZ^<?>4@R<PeZN>2WaX\Mea)-YX:+RE\(aJXQ9+,RV)BX7@W@IGN./M]aK2T+
<@DGL0-;[RP?UL<F7\90>>?0L^X4AS<KP[26(07JKGDWg+@5/DdUHL[c;_S0E,I7
-\2^#D_4:>:[7+eL(A,,c1([OZ;e.M^.^g;01dS2(dG_c:#TDSBO64TJQc)#Ub(_
G]C9]\#;<]JWEVFOOV,K6^&W)VP>94Y1F3>S-ECF.&MYH[ReJD.J]9^-J3A>+;IB
IW:cP-2E6NW^9731=XYTB]=b;WI.N>YS<L9^cM/U]ACW+;g3/1b@:F/)4AQTFJ_6
#W2;4,S+^AXWFYVb:)RRg<H8M93X)7P?]&aBc7>I#V?DK&:BHF?N2FSEQ_Q88WVb
IA,9V<4eBPNY,@7ceCX1(5#>R25Og?#WJ[EKJE/N+K\KZ4_,ZEPM\J>Z7(25V(P3
[,_5^LDXL5Z8,C_I3/gY/XgJa)Q@+CYKNQ:B3b/f:XZ@?U:WJ]:FQS&?;=f(XIfe
B86)EKLFT,31MZ[6K:Y5KS3gH8L<E=:-Z5?Z+KH[=#EAR?HL)7RMHICW\8GTN9D;
e\U3+Db0bF/dM&LCH^&E&?MY(4-0A<A+fY4D;GN&QA\M^9GY?.+6H0UYFaAJ?_5g
42_:TKIONd9a=_PA^-./Z+V\^.WQHW)GXb&H8H^RaC]0]4A6:+_K5(eL/;Y=I5[:
Udd7)1#-aF.DWWV5AdK8P3U@)LJf@?Xd7S&G_(SO[)G/A]K@6TOGgfK8^[NS)CbS
cXY/&GPRaA278gX#1bOPF>0-RVRF,>W<B2D#0?\Y;8_,\WfIU9NfM:_ZS[e4DE#b
7Q]YV_fMQ#7KA8@gV.QT?f,H&=LS<T28JX.LD65FE,,4(Q3<d4C_[ddP9//O+8g2
GFJP,c=VD@)N2Z(BeZ3D9=]Id-4UD+g;bX[:&V:6H2<5^O@PRLZP60Jf(-5/3GaU
E9U+>=Q9?FSGFa_M@RaUBV6S8Bb^Z8J/O&<@MMHKVcC[4FR1)d?=ZS#)@@gR:1gd
4V,Yd&QU2Q_fF+&-X/8YB8CBLZFK65OaY4G24+<>D29>a54d/M1&0N<e9KSBZB97
YgG\dDD=&SV<.UMRXZAA4a1IaIbS.aR@J&Lad93B05^8WSc4;JJ6ecM8\-gKGS=(
4CK)[4IQEU@D]SD6Z54@OEORgg=L2-d(\B5?4@18b>+SKc\Y1@ZGC/.2X/:+8g(F
g\T]cUgg1UU]3@958O@1:[13KL\I8Afc@A1>>(+S]cfZN-V6BU:F3/?bA:\[P(C8
[9U[OKJ;M:1C_LCd,[D>e+fH>13IP^67I59.L8aM992[(^&EI>f:#W/-M>+PCOO8
?_=Y+&DYPAe-F4bTe\@fZeP4(8=A5NJ>e.egb+?/2;0)1LML7@>)B?]?S8I#7<g:
YFJCZE&[b5)9fG=(Nb1Zc>TEfS.0\?-)\0)^^_:?dPH=6Y0MRgGG^H(^d@L@;U+@
6aLJ^0+CQK@68^X5=0Jg.H,W9HRU-.FQX[G6JM+^Y)CC[AX+3YY[NeKO4N<L:]8,
ZeD+&)62.bdI>(MP1QM0.O)5<0eGb8/eT@ZLGN,I\?])#a9-?a^A0-\5ZWO#EC?U
35LD/c(Pdb;c>>e[>]dAQAL;e5==[8[a0\1;:1f=P_VIZPJQ2-f[(FH@NDC^)?5W
QaBO<dWUD\e(,YcUUYQSLVP&Y.5[[BFNUGMWFXcQ;_WH[;b-CaAAf5&&bW\K(4D&
;@]^^AY3L>H\MK3K66G.12/?a6/Q:0@R-PL,&e/CZ5&=gI[X0Pab3P<_6XT(9UNQ
.>&6NH=F\1Sa73E)RQ<SLO;YD<,Ve\bQ\H7)@O:GZ&RB[]+52V;P#;PgR&/&;+Xf
@5KZG-N\CT1FH#OOO:f\CV48_P0>J^fY+7,JGAH01FTAU^X2-e?#H6421B8IO7fO
>0-LF+?1>F1&a&D^+X+,\V#]ENZ8CJQHb,VT(PBF3^C?1/QPT^.Y3YE),c_NM<,[
.9a0:R\g6b8D9)H23bM20L2E5-&5EX69@?Xb)bDXIBQ.M)AcD8#4bSTFH48ZT=eS
W^0-6b;1#H3aX9O]ZCJ9cBOECH\(T;>5Lb>^g@)//H[/OCL6FGf8acW44Qc\V_FK
JPG<#>)JX.VZKX3FO=?GXgM+c<EWE-#2&OV>=W>6N08DJa2F&D25#fb1_F\VZ\Ud
;U1QWG1?Q:J?KLIf0FaeAAW\@9XO<ST7RHf.;0TVeRMc7]GA;;X+30<[=-JPFU=U
a+,L&8Ra1==_?7(W:VL/Z36+8I(\914:^GH9I/cQ1Qd+_B@TL@Ndg#e2Sg6&PZ4<
_gJ&0a/=]B.]/MC_)OX>K3A4;?M5]N8F[R4cgbE^.)+;:;<B7.A0EHfJ^)7R4HR=
b#,e+V?7-W/;CWPZJO\7GM\-MM<OZ2(U9aP@PCbTP<#,-8\7MXKTF4S2:WI6C=#8
YCGNIP5FeYA/VH;H#XL4T#b.U9D<1aCHA@.I]L2MD5FJ:],0-F\EfU]Me9fSKgP9
4QV8dD(^(&(^;I]A&P78GbZ0]]-P&XF2?A/)UPfdReI7/PgH4X,2eO,ZHCY;K9DE
+LHAL7=)J]QbJEUJAf7RHU7-^/N5.OB#ARR&_\B@U8WbDIg-(XCe(;R42M7?P\3#
QYT-G?+gTPK=RPbd\4,VM&/?7Ree\d/4CV_WSf.=HS72)66NeORB<6.V8B5&?dXD
P(78aQ]L3:\+40Sa;7\&QC3U->NXCTBKJK6Z+f:MBTEM<G^;cY:\_NL1)&&J&@7=
(6=<ZFX_R8KOGCCC+W^EgM]G3ITV_FI(##EgR47EOO0MISRF>YW1Y)eWG-B8]E/c
=R@9>a>eR_#EQQ#DYU]aD-7=4,b-?P<]@+N2COAJX>F7AA7VA24QI,8+4cPAWcYb
3/_#GCFR^I\W3d9EP:<UIeP(6+\#70^M42G.&8?bd)&)W7/:[@8D3d-#4T0O=@fP
gN]L@LC5U<Y\3^:e,7ZfMI#;^7MZ09a/Pa;O>Hc2E:,O9d?&gO:2?)4)H6Lgc.ZJ
Q&XEg2(D/IXHK;F+8_C])E/@5L)O>NSH^6>=^^DBY;)E4g/XKK<+^PV=X<&X(^_)
^gTLe5>=0gg_X[[KIO]K@EF7B,PRK=d;#gU7\e<g]b=[6<)G1?FS887J6c\XUZ(_
;][RK9)F?C3H#RHdM,)SB9J#1_b3D)BA@FS<8,:5+8.:<M\-E<1A6&]0NV+KA0QE
8KP,L?XA3T8f-]ddHH6B5CFe6JK<-)+=_TZ(UJQ5Ab),3YNX30\9;M,gRKH_1L9+
]=Fa;4B):25.>eM>[/_g0XIV>4UdS.<e=V47=1H;ZACc3UQI,Ma9_E[c8Fg5b=2C
?gU84Lg1P@/B5M#X8V0>(SW->Yc\L(G^IWPW+5LCRT^XWc-;]FPE7PQZKJ30^FaJ
JR=<L;2E=.1_0?4N](SOUJ7eRDR#:WUZL<_\Y7RWOE;LMgD_ARVXF30?WWcB>Y-1
5.d.@&0UKMg931O^U:+AW_\dLH3HB_1A+951@)504E/BV(PKg8)>b:;/75R5\_62
D/UCS+Yb>?TT43R>#;,S@&93;]3(ILgSI>]_P84Z1/RQ:e&.M8S::bdPTOSL9[c?
]YQOM(T\<;-6cNM[f2H@/_YC23JAI>@<JV:;L<ObEOC8^98\#L]C3d>]2X=83+H(
X??2K<4KZ6SeBZXWad#?56EPC?\>?1(=5JH.2<V[(:<VeT9>N)C)KJ_eJ&de7WH2
Wed7/3R8b5.,0+=C\JS-.aQFV9g5)Wa/cb2UA+=,fEL<Xd>Z[-2BDA<A)f\IO(g+
O&C2UB:7_^fF+;;2K]Zf5H/->./f3:LXd.:9DDFLNN)NK0YX1/R\5^83R3ba0fL[
TF@G?eS3Z1]>,:8>+_D9Q+.MHO.4Uf3H6;V,M[?6JUL8Q)<0VYL8,F]L,-[PJ_3G
W2MFg/1:K\=MZBIE8S):(NTfCEcB6b(8#4+)VFFNT18TYMTZ\/cd+A\,bQaH(N>R
Z.gTK7I<G\P\S=I6+fgDM)ORU;f&3FS=f8//7R5#DU3GgQb22D-<d]+:>cBG4KOC
)V-#ZS,89eD=7d=5F.,R([/>eDQ8PaIG(N]/F&fPV;8\^.N@MbV:2IE7dKI.cZf@
Ba9&3-B1;_UWO13Na=UOKS\T,gfG3-;_\-O-.cU;5<9G#@8d6PUPRGEcd2-V7(c=
YSM[78cURI)^W3#@db6O08;5,R0S@3NO_Vf[Nb>:#U4H.Z,_<49/g2;].fM/.55;
]G0:P;b:AgY;]FZP#R2g5)f.e:=^87aB8_W2MS.?M0^=?@9ZU6>V#QA3F+0_78L&
NYH?J>?=:\7<68IRQ5I,Ig40fKX5,9USUZB1[b/W+N#-?^])AX,1f,JbD>6R>I;Z
;Y1e(f1<^N(M9+B3OM#2ae#CQZ^NVW-eTCQdR-C_14,=J]d?>JbZ^-XT7Kf@PYa)
A;./K=EP&eM:#9D+IK0.76^N7caad96T/R&Q8-&fP,^85^;UB5)3E=HfMW_;F]F(
T<A#)SfYGeaKgU3a)H5LE0_RP\b/REHdVMH5b#??cb_a&gOYU5NEYCDBfT4JbFg;
@g^/RaBH?KFP5d<5Wc>,K_[HZ^P=Z@DS@7a?^BOQ_\(NX]3=Q5.cPfTP=::/;G]e
58:#?2(@gFR^OCW5W1e5W[fSUc:a=(;ZGZXECcBABX,57CP=2FZ<JPND8c]ZLQ[e
,,X<N(V:e7TaC6D/d+bHS.+CY5-OSHd0RRNaa]ZdZM<5cSKE5(L3)W(09,)ZPZ(4
US,(+IL]Kc]SPWPCT]B?15,H)6SPRUOBHIM,U1@54Y:EUU=-UNBfK/EP>9cE)ZQe
7<LIL;e+R:ZaB.f4R\aaS8c&b.;=3<-6SHJGgI22Yd\<fJCAYYb/BL+EM<//Y.Ab
?RX)FN0E-7@dOG&Xf0Yb=e@C89Q4?+<;Q7MVJLN;Yg6:SF/D#Ee4-^USQ7\3/BC0
&->2RB4_D^;54N-<P1A-4DU9&a1(&fdW8@;JCEZ>]e9/=e8-;.e\&&(XBd@eb/2C
(:^^eWYIT2^3[>C3/,=2M__U5A@)LL_&a(<+ZW.W5R1T7AUI4R^+W;TC]fS?7)5&
FSDeFM5A&M?df_]&+(F>C6.LJLegEA<[5S:;e(]2PB0fRDY^.&E7IY\5cd\7T,NO
6-E+5>1g/8d\C6X58@_)IZRd)8._#4H]1NK]gEKM]4cfec,U-30UQO3)EbH?[S:N
-ZH;J=0bI3U5]KF1:/=V6O0UU#_MVE\C-#@]^a+G?I:R:EE9L&7;ST#b[+=:K=UA
#K_-;F\.Z7F;gVgMG9E5,I2)e3V;(7a<A<)-b@9YS/5847+ID&1V6<\1e&[:?^bQ
G@#?1M&cVPDPf2\XQ>4&a3M-?4-8[gRa;LYV+E5H]C@g>_-(H1]aV[@<J?]-6LM_
[@^;XXRPNM?dH(O^/9]]-3<d8FX>P\U^OfCgXCaQbWAgU\2(@8I@(..Q0F:N;[E,
=J^f((STOK?Bf]BDUI0cOZ@7\ZQ?&Q/^K5SQM;a54+4@.VA_,4dC3K@_;gV+QT+Z
<cQ+G)&f\8Ba3]737;>H8@3^=T5LNW)IHF3]G:Ibg06[9&<9FIP6S(\Dd0gN(3+P
[GAEH+H2Zg=U\cD7Y)-(2/BG=?39[T5[\\(IPc3VJ5D0NZ9e7bX_a&;VU8V,UL\N
SPK1OPa8^5EReJK#T<(GWB,AS3GE6Re/U#]eQ7=MXLE?#;(T;Ia6WCW,e]d-DP-3
-M.dd48IOOCS?b68KV8ZODHZ]H=V8MHI3?EVR8?/Qf/F^a_cd-&AYVD0L;ZKa7&8
@aL5_fVWb]5=BB.X.M&Bc0<V^cZV]+.6S)CYA^W/8T5U@KJ390+0Y)6AQb5;W#F&
(;;1Te6?@cV#B^,QGG_?cL,?cY0?J/WfOSBTQ+_]M=2?]5cD7e5b(<TK@E9aUY-W
+J<64ZG^WABRO6TV\OE,;E<e,QI8OfQVKBRWVM7)HWL[NWTaTYg^^UEP,>W2Q-9;
Xf;BO._OFZ3NH@;E1UKZ7g[gCJ_]#Qf409,&XWc55fLXdGD0MFgSD?Z)5TD&7C4d
eZMK<a](1B2db93I>IR_a^L+J&Q@ZfBX?g/&CR(IDOQLTB?AH0c]\:D7<Ff8[KX+
]UZGa>TGR>KYCa3(9B^UF4cfU_DAgH5_1)0IDe#YLK8?;(;Q-;)3DbR1\gTX_\YP
A\YW)eNG_)G7b&,W8_P_F;a/W;]G][V^1ZX\N,_d1I;;;I?X=89ZJ]I?QVL=^fY.
]L1-T&a&1M;>3@DMf,ZeKVJC#bIgWD6Z508+aW3a)-?KZ7E(]>T#<MU?,#XT6RXB
gcWMa2e.DN67)#:M<<WZcL8?gH-L@<A&_,AIK9J#U-LM(U<>TBK(OE+<ZL/(Zb(E
N,bWN5eY1RLcLIM<PM)Fc0;1_/3EED5CVM:=dFPeE:MP^FG3W\#9KX0QO/4&48H&
SHTDUH51>EcZY;K@W)2b#@A;2KTD(R7IT[P5?[VQ\d^IUP7EB,d)Qg(T7L(K9]&<
Q=&g(@[0TE#bE@_=T\eWCfIL+08.PW40\_U:dW[\IMc=X@d0(9W5)W^PH=HAZAV;
O1?aRJ;Gf2XLM4NGIK-JaHaIV(]O<SEK7X3_bRFY8J]N=,T4g#,YF6SZ2H.(DADR
K_PHBSdYMV<+U.eKDd,-[3-A_,Xd(.<6aZ#@TfYN#L&?<X0M+f?=BW/96e.373_W
V,I9[R<2C)B-1XUdc^G/;K-8UVN_-[&eF1P9dYAOCNE)\4SH[?<[LF\PKFT3<9Nd
O;;+_eSLZGJV43.7:M;fOL+#2G5cf?NY0WOWU8ae)HOD^-5F;8QC,,5Z5J6(]V?X
baYReB?0[K>+J2Y_9d75<D?A]QD3:ZPJ]]@L.43V;XeYK814?+Y,g^O&5,Fef,NQ
\YRgB9(,2.#U]a\TG[DgUN([.]7(^Q[U4YaZYS\1.FCQ8Vc)TU--\K0DeTA)A^(V
<U=UWOe_<?:8e?P<KM@e:AW+ZcK.+:V5(9NJRa^7TG5b6,^TC#LIVbf&S#<#;P[F
HQ#8/IOIOG_@&U0J&]W32<L1QEBE\N4C&@_^bNQ_]66\fCDeG:0dad>0B#=UO-KR
)C>6Z-ZLO-;JT-38=H86,?7,,,e?#W[KZQ;YRKV?AAP35V4P)ZWD14#-f,?>WD\7
KX&ddIYNJd+8\@:K^4>\,gD_:-]>ScZ;2]3STJ/I7[8]JB5:1;[#(,KT):UY:1>+
)9Wc4NP7H9S5JUI4?K6R/>&&F+f4fDXFWNIQ#B,d\>_JLFe7fcd._HK@Je0-N+D=
>9\15#4M\a4:[a@9_]F31BdgXH.G_JTa3((4[39>TB#-[FZ;@GZ-XeN96>I]c6PZ
,Zd+ge4:[:H,D2186UF-WE22g4WZE)/5_e9L@bF_>0>A&)\A7.F<YUJgJdOaKM3@
(_eSe+;BWd7e4NQ4P2g;3eaN<@;H4GVXMB+(P97MEA\HK>DN^D4&:<b,3Lf4;96X
(2#H:,MeEBDX2V^bIFI?ZLG+L@01>BUb3[^]0GWY[6Y7\fST/5agYN[Vg)Z;8fQa
O:5;7S/NAU=)AI3MG3O<>Bd.#NRMV>4=HB9YOPERJ>Df)QN#c;J:>;<=C1:?WMX-
GK@J>BFS^IFN?fJ]5Xd/_G<_;\KB:5Y@/?W-40=M0Le@dDL74<_AHDYX^I60RWDZ
N_QYP^6M;6.63Gb/0F9bA;b>S_T8B1.[e.C6VcE7709GR[D>3X;:YT+8.>DB]NX1
/+GNGT\C=-VY.FeY3^L81TE;Z2Y_7T.6aJ49&(gaY:P<JGfZ^6UK-<=g;@L7bY;7
RL-?Ze23b178/J1\E5DZ^fa#52]QWfAS:+@(M;TITbJS:[bA-:/E^A8+>>:&A,^D
U=YE#U\P^(.7)YYSMM4NO;&A/cK.+RFUJgL:8B9>J4W/G7a5I=R&LXW7N<-3@M_O
)94\5dCE[HIHCV/P#FMb[ZUd^Q435](9c:,/2<5b&6U.P:61&?3Q7.W/74:;c+^7
W>?-1MI/(g+M747E8F-[c=FeSfEB/0.(R9INQ<61::[<YXS-2:T52/P&cMRQ@>U+
8fH(#3]W8dI1UCRB3IV0IJ.bbgS=)aS[6Tg0N5A-YG.^H)e;E=#Q[,&bBa9NBdEI
/:V2W?OMTFE]2U&LRZ/9V9+M:O:;,gYc2g:4T\JB+[M9]<T-+;JS8c0Z.C1a?A9#
K>=ZJ&,ZT-N93NZ(QEG123+_BKa]88([5b@YIQ^6YYE^LZ8RcaXX)WNg.QZe[=6]
)&Z8Z]gCZ;V=J#X</KO,;6/cAF6VI>)a^GT90d5S^aJa6@4b(3a8QZ#RD_#,Yb]5
=N[-,32F[gZBO:LOTaU24UW:K6D.7=R6L+F\(<a<^3eTbP:/9e2PK&#D+JMBFg\:
Q<6=?gD/JaZ),#9=;QX1]4@:5TU5,5#)TKXIg:OKD3g863^3TZcH_34d@7@fC#<]
I6E4>PQRHHTb][LAfPWDX-gD^X&^dOP+^Je2dRK0M<H#2Ic<ZbfU.bOgfaCL#GXS
2U&28<[H?2+.6N3g&)1H5]3V@;SL]Wd7Sa^(Xa:ZH>Xe&^G^#0e1A#dSBAV5g3M=
(J,M/J))I:V04#@b84FfL1JGQ4KeZc)3-O-&FX.&33@a&VZg+G<IM=O>3U<4LXVQ
2Y1OU;TW7GHHU@\ALY?L03aBC&V\\U/(?aJZAJ]^4GYdW;P)(a)ECFV,#1=<CM\Y
DYUgDacGO:Qe6ga06T0@b&0SOWf\S0)F_#L#^^[LE8YVPcU[75c+-:9_V/1:<]\@
4<3=ZQAO6EK_bXea:H16\K62?)SeID2bJ_bbD[aZYF9^PD(UTTKUaFH<.5>baY?X
<)bB)-8,,fd-7+Yb:;8A+-&_fE@9GK:1@T,Q5,)d78K6a@?aWZ4PB&OWUI?Zcd5:
XMCeKbE/P/,X(EcC;+@B?4D.2RF3^;S/fNI;[J5?CL>2<N5<U.aHU-=IF>LggA_E
J6J0/P-<#065,.1/\&W7#Wf^L&AJ98/K[]JbE)+\M?:gL2?I&S(2[0A4L8NPU2X9
D(U4M>A+Y#f79;9eeE^.#IPdW6MHY#/II;TdGFG#IAIf,M55FG33+>/:[W&1Ta@R
N7<7U))#1W-X(d9-Y50]6Z7\HbTA0R^<#eK6aQ+f?W2d9_Y=LgH=+7E4.Sf-_VY3
@CRXI>cN#eHAAUbCfc8:&JIYA24^G@88BYMNe85V6QJBQ]8+G/5RG=L5G5U3f6R]
HgKcT,?CcAK80&A>@a29d:9.I;ZG:YFCE;Tg6R6cGJHH3]OR;[a:H/QE(O68/-+E
T9A_BXWWVP1DXe/[<4a=@&M6NL+_:X5Mc+&1]U>=I8c2W]6F/f-#dQP2=4GdFKgR
#4FQb_]M<TNf7QOUg7^[LgMAK9-JIeGAMK4_O^<e_T&C)D0,H;:6>P</fLVa#N=E
8(^ST?62X0K3:]TSO9VdYW>,fJG/5N-(4)G.HC9V#A_A6TI+3Vc<aK3UQT+/-\:-
.D7\Xg]@.e_a(_/F#b38B?XC@LTT)ZI5(.DZ..?[4RQ743H[5S))d^(L8Uc)B3J2
9N)3U+)O@=TI_=e#Z;4IcGI1I5[]Z5ICQBb^^QS;^,<&D>?_8b;-]\.6+M)ZT[H_
b_F(UMQ6EGCY,/]0E:0(0\d1LQF<MMO@6K^0M]f3/]@<aZ\b1Y7VEC8ER+<E0T>c
^@Bd[OK77cL]:W7?Y=4Sa#4f\)[7bW5W;4,R]YAKQ87RF-:W<_De_6S-eAc4JM0.
IUfCWO8@+1^5A&3G[5_1=:Z^2c,WSe3<F>B+JdKg\PV_Cfc;2_/Ub#P)D\Z376g=
+=Q?&WAgbfeX<[,:RZUW1ddAV9L;,.),JDB_SN+@fMO0757Y.+GWLX4/E&;GDE8G
S&-&bI#@ee5:b</b=30W[[]APJ6W^(c[\?Q+_.-QOEH[&)&b0,+/3eD9gIdKJ-BK
)59e<2ZOIE=-&g##9<IZ>91a)ZJ<5LD?R6]F3C_<Q4GS_^0[&7U6RJ>;XdS]eJ+e
H,g_;+PL)Y9(CZICPBL7MU@2+fBERXK/:6[2\IT<dDAT@f?\KeAQO<,;8F6L#;UL
Wg5QU\SSJEM;Mc4TSNOeeNP+[78P&A<P&9D?[ggD1@a=V&,PfV@L9YP+.g,?&TLL
X(+fI>Cg-/@9RY[g3FX+^_1V5@?H)[0/BHO_44R_eY;@aJfc__:.V:FU,Tc+18PX
\V?ag0/-&:7<D/dMQN]FB-Vb?6NI]+SgOZ3JP#8R]/.0D8HY1KJ&&7(XacD1.62:
fQ\.Zdffd_AaRG_0\HCeV5;NfMJCSP8NW18f1L)Kd11LDLMMSAK\&[gE&J+9H1<_
+ED1+NR-FeU_)P:IZYSGW(I(0aD4Hb;U4e;1O[-F=2TV+,=[bb,gZ6WS,@M5_N1O
CZ:W:dU2GZa+Nf4IBMX:E<X\dKXYSYB\?=AT2D<bUe82Hcf+UdCIC;c89c@[cMU_
[6aW8Re,2Y,ODd-ES0BM0A8F22<Q+BXR)7>C&0Y[-D@X)Pf#]CY-V@6>\NA612C3
-CaE7TeX)\B1fKbJ4S,2Fg6]<,#F>d\]U96I>a96RXMTB;bIb#g#[fV:RURWVZ0g
KP4U.ZGNULR^gH668fBJSE5?FH0ZL8,:XS&fY2,0<Kd4Cefaa+_FLZTTO#]A6]3.
1Jd-7G&8SdT+@O<9+/[L0NU_eW3_P^/GVa)3WeZHB6+=0PVH?_A5>:,SRVCe6_?P
b8,45?1Pf7aETa=B-2ENIM>KcN;RKcBHbP@T20G4Ta=cI.<LHJ?P39-G>]:;EBAT
4+gM/41YX8W3;BA1+,c^9G:9eRC]O^)E>Ag@dW(8=OL0/b\=P=D0Jf0OYWM^5)C?
Ea>6<Q436S0OKW;g+b&0cEKTO57bbTNL2>FWUH0OO)<^U&8Z_bfJc)cVPF0d?Z@a
FU#.cU]KY57Z=G[?5Q<#\aETgF94<PC#c+g:+]\+TP/f:BX(>f/X3G3I\8g)Bf8=
C79G0dVZ9ID+9J<TY;>eI+Gd?K\_1),b-G]AKPT=CA3d8S_3):&\gNS<L.3;;3&Y
fKBK,Hd<]Q#Z\aDKc<cTMFF=14aQSSg;F)UJ+;2bWI.e,OJVP>D[,_d).S^U;;\4
PMC4:@I2>2D:BU.c6:LR9eD[F[)aM)09STW8e&RH?S87&4P@7)AHfW4;&EGFW0Bc
-?F5dfZceCC0MS&<b0[(-BN=&QW3O]-O[2?0TgQHFW.b@]_<87+_@V]N?,3UTH5;
1?,X7:f\]<X,(0bAg-HCRg:,:KK;=gQcTaeYB_-)[F@c^:4UNSc0:M&<UcWKA4S#
]MY9c,6Y>bAGXG(.U6)^EaCM&#+^MYb1R[cgSUW4ZOZ_O=\+8eQ&)ZMY7X+/XI=c
1UfC?E4X29S]WX(a3VXG0RF67a)a83Q@7fRg#30>CQ(db-=Q3+?AQ-8<MfM/e2()
;JZ2BG4Q<RNWD_BL-)E(c#?;P?L5a<10:,:4<1[YcNTS_<=CP1>^G.LXcD\_V?-:
)Z_R[XA.VTTU\_=NJ&]g#Q(<.Z^T-V^bW3-8^7?g.3.JC\5D]7STP.;W/eN-S,FB
M4PSH44SQb04FH94eBAdMQ;,BCJ62\C1KP<+?T@U>eR0^g_dgV-B8d3D<^_A7CB-
Q\MYef:UZ.E/6YZb,@DV.f>=3,+f>,fW^2+G?L+X\I6&YVdMH=gI1BC@&+5BKg]:
=Ob/XM>(<IQF?a-G[4,(U?7N?-S/N?f[P>SPSXH0+T1?@NVLYO]dGR34>PPU_[52
SGA)5>J4@=JP@#>3=902de?.QEN1+T]T^W@+DO;L0M.F(BLg7E9SXdb]VY<dR@?R
?-/dbA@gd=J]UZF^a?3)\HY.B;[-&=K[JXa&<JIX@/,d]O4UJb@_TLLd-LdH4,<W
)cS)/1&Z(F39COLD<:X=?@H>Q#.++;Z9)CG1c4=_c3TWU8B7MHB:>\XS+QQ;HEE&
5c561a=^^NG;(6>O@P(9MMDR<_K9]CECO);eHOQ^Be[De;QD29^LDDG:^_UODB\Q
?IK=AD_J>GA?O;4+AJ0]d+9U^6V&=EdD;BJ^^7-,7TQMJGI6c5=[,KTLNN):?B:S
R;-DGYcIdSTc<^SA=&-KALJ?YX8G:1Z]f:aS7K@3UBaOIdO9Id,]A,fcQ:5[XAGV
^U._A:]-BKb1G8OYfeY]3O.3O;@[-aOHC]Z1YOHJ@R[XRO47(4/Rgf(#(Ze7YNVS
H6YG7BA\3?E.JSLJ@_WKDM2aWbKGTe<2T6831-@G5g&Qe@O?=IT;9.Q^6B/K8ZDe
cEK;^f8a?M45@)V\S&(@#?M);>)K5O#D,VbPL9+&,5UgJ=.9cUbfKTRRMCZH9_EL
OS2gJ9@L@3R&(F[AL0P0V,&XLcOb]Z(31)E:L#V1W[ZCg>5W]aedRN;KYDL_\M@.
FQ/8c6?60KD,.c_0=D>;1X_KbQ^4,eg)D&K0U/6ENAZLI.ZUE9gXR2X?\1/^?EcM
XS&BK+U(KgJU?=,HFEC_./:fFCM:U-LGgL:V8BGK0a;I510NPQ)\3A\8GN5C/CW=
&<-[UP&4B.1+=P5OV59#:\V>AXIWC/(H587<_?VYZ_eZI[fdZAD^9;C8fgC[4E@W
3#DZ,a?N42XRL:+KU0578[5f48,@Y<4/:HO.cR_X[BR3/eZ4a?V0]8]IH7)5[5,]
(4c?MU>RX0F_gKd?B?O0.CaJH8EHEKL.6[)ISV_LZOI?X68ZIA<Z=)cfg@<TMX8I
@UT8NTf(_<YPMY+H4+L<^cHe)2ZIOeWQ;42/c\],f4MCK^C-W#J-0>-B([&);/+T
HQ1Z3a0?6/ZWFEaCT#@I@eQ^f@7+<Sfb3F(dL(=_2AYcd\=.&,-^&4-NfQ.(XVU@
bYR3_b13Z]2G<FLPVU2E[T#gdF2deBDQCfX=f\06ZZW,XF75N\dU(/-E:9WBK+O>
JM[XK51:XOR8T=PR7=P[1D_b9-bST=/:3#3(<()c.,[];W?F)D6ZO]c]5961@V9A
+^=M@aG&\>+:KBUY>KU4-W<Y+Cd+J>R3H-.T3/]M4L9ERPQWY6YQ4ZRgL]O\ABa2
_>-7b;KLMA=BUPH4Z<?QI?,U-6;HI.I=2)dD=D/WR3_#\Tb)A6L(#d]3Ze&_JD.V
aC2Q-L;@06Z150Rf(#K;TcFF.PATD:]VUP\H>eMcg2GXG)-X&d)I&?98B+I9:BG/
,KX]?R.[UGAe9DA=<GC4LO5a)>6HAC7geEHD;K7QS9YY^K9R28.AR)?\U+V7LFP2
a/E/FLX#VS@D-)f6QcXH[G7[\g<Kb@&TO19RL#46RA#fUAQV@\;K2JS13ML#N_3C
+Ze</f[QeMXV&T5N0cG-55cC93YZ0.XE_)A)FeE(/A,&&.SAXQR1dUYHg:Lg2dQM
a#VeL:gPd1SG8ZN#JI?IcY7FQ8bOEYX9Y:?J?Y&[09[XM<?:K=@RP[f3R(HFA;\#
F4RJ0M\.IP&WD;LQR2(RUXcc\ed0eFY4b8I72+[73L#af1)f,N+N/IIfVK4P>+fS
O5-acA6e[Ya?&U^#HDXE8IH0LKcYeQaaVMOgW)URB+]0deE>\PE#U8?QT#]O9>B[
eGE@4EA9ead_+XCA=-3_K22#(0JP5g-+AUO\/R2MB5C.E0Rb\Y2E,+N,2gQ.3A6=
62:,L[5Q,dL3c5R@@UdH/-Y93A)F;PWV4[G4,S1?<<_5.0Bf1(#GHFZXL2C80JWG
a.B)T.#<LcXN1^E(e5@6U?K1C)0bg<9FQ_U>5OX&WUMg2<@F\GB084HP-)f#C.@6
BSKd.e)4X<>>X[>+707W.=@)Z)EMXW]E#Og\[YLVW>OY:#/)N1_/EIJ?SS^V<1J7
?D=IU),[3PI4aLR@8::V00b3Q>4&#MEW3BU;>N]MN[DP:M[S?&[:J:8F5EBCE\a&
B?)GMMB1(D:8BV\P#a?;LabJC<bBCVDf-&HW&dH-7,If([\OQ[deNag5aA7307B=
N(;R3-VHSO^d>K8G7NA(QW@&TaF->NOPR@..O62:=WE]D3\#(NJ+2a.A9VO6#d\3
7>AdWNUc,9PY<[M/1:\B]BL7/9G>I33>:GH01UaDC8eLEa?=;QP]PE:(MG(SER;Z
-e[[<eOE32=a=]M+[:R(Gf4(,\NVE-R7//dY4(GH..dD_1G>.A>TYeUD,E+Gb+gA
;O7-&?60\@T#(BO;)56PM2Y):-fP<O8f\.B-.]LUO2?-GW:?5#a?L?157^=f(d]S
GFY8EDELXDA#0LS?0SQ,+gb_3)4gI#..faFMBPVYbR-4W>0@N-g0P^5K2(&1QG/7
c&DdGIG(I(g^V,ab1Ve?M76eI;Ye,S+[aK]5PMJLTJ#;Q4aC<g?:7X&EQ/93/-g,
4?.LRM;=<6RSY):_,,OMQ=A2NN7=#(=>NYU/&aMZ@4W(Id[276)I09>@V2G7V9IX
L7035[Ze@6Q&&TVI^d/N=)=cATeF[WUEPPU-a8V5Z-W=O5W:FO+D5:<b<eaG]:FY
FR&]W]e8XX,f9=4R]bf>/ee4V2&C#\S=B_@bB,@+McbZf7__2WMR0][L=<#V5cf>
8@Pb;-9DeFe7./CEKEMY,LK(==gaZK_OT7\<0D<+f1gZ@SW47?OEKL-:X:Oeb?YJ
/&\7cA#I,PPP;C784b)MB/N:)fF22HZY:d0fdK?S>NA=N=SB2<.Q9gGJWMS\JA+\
2CO[8.14D94Q&>9/=V6EM5>O-#0LW[],45(&:c@O;f&V#[3NM_?QA>XNbW9Q-#Zf
0N<Y-[H,4ffg?-4YF;;7aF[ZM.N==>:LQWLBd+4/RYeY.ONA((,c2[39V:-/02gA
&S-3-8@<TA)I0+D3OZa5YI+G^IR1-^2=/04G+aUaV<#BFg/^T+G9U_[_3C8BJ4(O
3Y_E#8<P+G<@.3/(N41>U@X03UBQRXBUV8<a>-++W)+]GJ9&8[E_WN@7.:>RBE@;
dgL>]f>ON/eF&2A6W6M@EQTE\]dcg^N.GXB55AI02-)D.]QM]]?T35F@V.8]LQ7a
H=b;4O+f#U>bHa0OJ9)>Jc>ET.(9Y-6(0Z_[(>58-AA&.GY@]1dQ@Ag9-c_Z7-_-
<0;:=,V5]Z]#(#,J5)VK/C]8]#G?BdNTS=C4LH[D&FE?DX1)F];-)c6:)7@&aBc)
5&&Z6FG/[,M46fMYF-O\[4)B,509UDRUU,gZ_9-60&QZ/6S#Pf[>Nf:4#8a^cdNQ
cU(HeLNIb-<\Bb,8KUFCR#=Jd:T:<0XDe:,P<@Z8R1gAA.b7?T(BE7O-b\P>YbGd
K-4>JNR.YMSb0OTDWM5INL.Ob\S\Ae@b6:AYQ^GG0[?1WMUP[I(#.^M,6[/(9BLW
_:D2aEI,F]6>5#e-E(f4?&1CXOAHOeE4M;gJD=U0XW]8YK<3OE9FMET,&9dJ4VC,
A6?c4+J&:)]CHO5(3K/N2Ke?+aD-cX@CD]#0_AO.^9OLP@,gH=.fP)Y,QMbK=dVc
aFWcRIT2V]J/:.V^eFgUAPL=^T3LB/_7=?b>0U]5T087=<BHU(1YOFJ7@L<73JV-
YWA+^AF:[(\V:<B9REL8YOQDFU@@Y/a2<b(J.6]a]8T#:^gLda[A^P4^5D]f/8C1
VDWI1=bO37]eDYd(CY.5>59X27-=WX9bG5GOC0J70GKe_I9-e&6e@,X@BK]1NeCd
)WT^bKCL9eJH1&6N^LLg39-f+_.d3c&Z/@RP(:+a6;H1MA))g7E7;a@=H+4Z5Pf\
#GP=50/L+@7e1D+O]JZSH,N>2K:De@J6:=Z3#a6<faU37).1=-_AZQ)@C:IH1U=;
\B+:;(T[-\9SN,bVX?-],^),M^,dJI62PQ<WZC6.U][O.Dea)b5-Xd?5Y=JLE6\L
QQ2a#N_9T/>Uaa+P+NbN>)bG\1]P1C@3gHQ?3_:H-A<d:,RH:OgL3dUX\UBG1])f
9>fWgS+@8N9&PH8,=JP#b<0VfB[+g1^B:\F6\J?S.dRYWE8R)H(?ZGO+?7Xbg4(L
4O>T6CEa184VF5Q@CdM=,3b+_B3-;(7>UC)NC_EE]bYY1R;52&-&930\I9QDQ;5[
#V6NP#P9U[eBBGaP:#X9g)a@-,H,5Ia#OS9OUF)a,2N3f3Wc<;-FLME))gUT\07G
M2V)],.@O=IEV2g0Q2J3Q#6K_(7NAD9OP1AFGXG2;NI#0?:e2_HH@?S\5NTcPHXK
0ZBe^/),:NZRb#M=9&B?N^2&g,HL?^ZOEYU;:UNO5V[6J&N[deW47@-FdQO-H#8d
XLM<6TXJL>aJJb\eTPUbCc84-9U5HYXZAN]FZ7;8HUe1=gBdQEC>[UYX(2TPWX/e
<(+eeFb]:AQU6-\e#<A^)0BNNPWMd4&CJT?^>>SQ760T_@=^D-M8e+#28\(IL5Y6
D3K\V3PT.a#GWARCF3Q;>8;C\TX,=If7R[)[^7LW1QO,\X>W]PS_?,8<IK\M95GG
OKVI-SZU84?HWGEO#UDfeN9.9b?6ZTbeX9G\5P7<]JMBT/Z?:SMP6Y-W35).=P,Q
)IJ.+V?7Y5:b#Z;@<-W4+.X,dX5,.S5#=9.#L_/2+L55?d]DC8G;TS;(/>D06dab
)_JA7Z4I1V_9JU7:4gcEOK,C8LLf,0XKI(DT>VGU8=_bIgV:6XIB_-EFBUDcAX<F
-))N[T?YWY)aCD-KT_->FLGC(D]7F5+#Ec:2^D]T]H9(:XacdN/1>VP;d4K2]\f.
KAWUdbL>YBC=8[:1E\)\V^CUT#UE]G?B3T9g1,__+c9cI8_#e)KaXgIUDaVGGH,L
@Be3c9XJ(E=Q6QD_I\K5PbY&>I76fd#4Tf\f0AF,_F\9I(ZYGB^K2=NN?1-0e@+Q
J,SQJ-(3-)TJe#-SV\c_>WK3<RZMT]cK-M])O#>T62g\JHfZ2GT_5HFCWRC4(cB?
K<f_9NO64.af\9=fAf;FQ/Y\ff=R3>e(gXQIUdSYF:.dBMAC^F()B&L,,Y[JR])=
-L5^4I>VfR#DX+2^6=e47N(gW3faaPS]PI_/<f5U<3a^.8QB0QHG(fdX4)5a.(V<
/d\]Z]GX;9I&<g3)58fNG1ZUZQ4J_@0Q.<Z_;Q3Z1M/aOg1?MX3008f&Sg>QJg\<
DUU.T>^67V&_NHeL#d[K1eKY_[D(V/@47;a(UJUgRPH/fG_OeN>G@8[f@&&SQPb<
W7SGUD0VI,0F9\JQRd?E0_8VE,Q#2>WEe,c,;HCHQZP]/XU/8[:-L^VFZW>_SFLY
#aPNWEK5\(8a[g<)bE5V9_6,5E\[=5Q_-;S&18@&5fJ0H,JKaCO=J;KMC\g=<6J,
HR2C?JW[XVK?&O0-ePZ>AdZT7g.YdZI12LYI,bR]#H[A0/-0>e<CT6+ZI?SVF1A5
dG+)&+D)KH.(gM<+:/8c:9(@)VP7\LAY91/e5[SEZGP:\0HM5;F77e)gSH1NIY:&
63&.f=2C43+34W^&_V3/J1?EcD#,5MJX]fb/;)(R69&SYf+]5gHBMZ/LBBeYb.2N
))#?[3;;KI3bZB^[TNZ6;.?RE#F05ULCeC&T8JVHIYf23PbDKN)Z3Ib;N)E(K5^0
0O(W&C<Y090d6PScGJCR@A1([H4LDb2EK@=7ObNWTWeV+X(Z_FA#A@F?8b:9U95C
#c@K9,=P-)7.FQQ9F-)A]\gZ#DNcW?c&Ugg(WDO1/0e3b73cf-(2)P-D6R.=_@V6
8<+#VNNWB+Ugf>88/_g;KF\IZ.MF:3JS=^/4^&]HJf.>(Ve20P=P758G1a[FRN[6
FbR\#ZCa=&<J&KJBI5]FT(K;<T1LQ6X^a1=Z^WJg0K2-X;BaWQ8gEI<gM:<f^,NY
^>VKJI(Jfe\:WS1L\bJSZW)<\L29]<WF@#PZ5M.LLGa6@YW1KV829IA;)/UMU6VU
2>/FAfcQJ(KZS,eTB-dG780PPLF^7:f.#]V#4gV/(EV;6SK^O;_:+18Y&0POO3/2
6gH@dB@:9LGX4(&Ee-I(KK:>T04f7U)K0>d))E,9;bW86H791Td_0LP)f#TBUUa:
Gbgf;J_WY75FW2:bQH(GQ58G8.;;Bd0(MIT#ZFX<.]300HfX?Q#:NJ_dS-M/NYVP
^,IdB41JT1#VE#Wd1JL&F&L]&B]12R4>]I1OIKU,DA,_L]^+?_8RPJDR>Z3+U@7Y
4Y>fB40EC^/=-XYU#/bJY,X1G<(E(6]3??g.:NNRLVKGD[7WfTDC[[+&O_?/6#U_
DcFGK3fUUY_We]<V-+UGAAfeN#48QSKP<d?aX64(cV=_-SI=VHP,=J6JSU6(NbFb
-,L,-<2LO27bdNQN2P1#X3\9#RZQbM/EEg)+5CaAUR#Q,?K];4_<JR,0FWRR.=S8
XgWM4f:@RQ=a#ZIGY,3@;5HYKWPSW;K+-C/L<,XKU7;/f+g1]D_ATRZdS&T<E_\G
OQIRGRLM8@U/G^T&S(G-?22F)NKYE=b8T-EYCeNEB)T8=XK49\K@[?;?FY_41/^]
\Z@]e3X_X5aY<g-N68e0639;:\G]X6_d)DN/g)P1aXMK6J[cA[:f,/168b5-I3]A
Y&C>42WS(L+T3H(WX-<9DFDFc)+;WF2E>fgD;,dMVA=.ZI8Fa_cKf4RL#HVMI#R?
6ECeL>Vb4<<N\@gS?5L2FR6P3X1#9;/F;DHNc>&gMLH<S-YP/)BYWEWMbDgISEX[
\faXLF3S\1@5IHI@EBVH2-W&>BB,3,GRKN@((@25J;(<2[[18C_,1WS7B+-0X\6e
X3\BKV)5Q6JG6YY<67;?U\6_@8->MVF0-4:a?H#5EZG8?8^\fG=[@KJ(ZE;Y(KDX
<][.:FP7AE0(-WC5-@+/IC@/gce1+B;-1:=B42T6T5AB??.YRAL][>2TZVF4Ba6b
5F\NG;(/F(E<ZNb;9TV/c72?@4:3NFfa>Nb5_#XQ62/MYF6E.@ME]K&^+D^[^J,a
6&1Z:66\eYJ>gKd>^L()=,G1a1V,P.=_CADe_B_@(WQ7-_/fa_7dSbI0)W^AV]D#
a>K-3-,F:CAAggb;R2>(FZ;eSNb9CJMPDP4TO^T/:a<)&^-Rg0a(EH9G]=]]c#Ef
f5#P?GL=^J]eOM4WVM7Q#X2XN),/XA5ZMcAOf&.@<-4WZIUK:;_5F(NO]c2K402&
_[RI7ZYU[I@+(C3P9b[&>G-TOC/a0cS#&6]LT0]a;,^0RF\]=X)Z):DFT,9R)E,D
>dg;J?=FBP(ACEV=QH)>;T[3D#Uf_7Y)A+#/MbHR,&]QNV+(++A[RIY]TEVeKT0&
+U9>CO4;-D92a.329e^BMe+b<d-:(K0e]4\W(WeRN-6c/F82N\5C3MEAb+]>29cR
=O&e5ZQ,VC8.g<&/)c8/(#47,TF,_S/[cU5?-<bcN=Z6YHGg2/0^]H[_4JN(_YBQ
@WP@cg.AD9^[&&T@>6IQI#I+.=g943gd<FCRCK>R\a&Q-8NRQ[+G+:B.(EHa.<Da
W<--79K;G;ML641ad>bB<7;&aIPIA96fAS)@,:OI+=LR.OW@XedP9_P;,\&-YH8C
FQbT]c\d0Y+;>@]gT[W>47A)E?Z[)M^]08Ze6O=.=NK6MBe48A.SKTcI[7RL7E]D
aKeC9V+XKF4g[UMO>T,07T?54KOBQ)_:Hd#FDJD6g3&<E((GX.)dQD_:X6Gc3<Tb
.0^A7&;5Bf7+CW-g(KNJ--=2-TP](=gQ-GSKd]Fb+aI1&65[J83&8@AfU<eLH1+S
5@1OVH]-KL.(_L^0\I5+&bWBS5JaU]>-8A(A8#Vbc/)RY9)5#?OaS+50a+[UNQ&3
)9RNBFV+CV.O\_=309FE/J7P,]S+/U3d6;Hg772_5>UQDf8LW)/U#QC]f,9(+8>d
^[+SS:d]\;FV<cBODG;aV#9]<H5d[WBGgV].M(_@ccRIaDBTUL.:_D@6gJK.LVe7
4<[<[>-dC/BYc-W2JBGFB;)3U?(W^^_g\FO3a_4,AR@?BV3K_6/:9R5dTf1e,^-<
Oa.WGI&9GISPQ^c?ML/EI5UTDUg0:?DbN)5.ACfGIN#;O9]e;HYc,;f0]a:W;7e;
QD=2SURa?g,2fc4=Va=Q-IRLdZOHY#R3Y&)aGfZX;,U<Wc];2d=WNTeY+)gP?53M
_V3U3P7ZTP\d-&?#_</AXcMNdQAB_b+[\@E_@48g8ZAUeKeV(F2P)QOCb)J2O04#
@^=KFA3W(N,],,Z7Q,:D3.2^V\BG4]NHc&a+&LJN@4V<1>Hd-:S/\9E_UgR_cId_
T8/E?WS30],^^c6g1)@LOa][W5/O+aN\_?V3W1E@0T]];L2;WZ(5C(1_gUHJ9Z90
<CYV_/W>,.VY86XME?^Z46Fb]/-gLGJB1TTA2(T[V1?T_N^;a26f^-:)75b\H</d
1QI3E(+YQc8LI7GPHDeH[@CdHLWdfG++RDE+f?6J)7-DD=PZ[:E:R&<bV8KBXW9D
?-;=#&6:0b@#RDBaA[;F#,LZW@8<+^@NRbRA5G=-f9.7U<T5^3fXS_GaTPb:WYAd
?D1;c@&/^<51GL)[KfF19V@QaAP-=g204e)9\2^GUV:O25JQSfgK<_2>8Q=//&gM
5SVbdcU&T)d:IN68FWRAFHY59Ya,bA.HHK,MJX=eM^Y2cSfN>T9>;6]7fY[_5(,7
E:0^VDNGL/<6=U6G[@WP#fX\Y,;HI-;)aM)Qg-ED?6Rb<1c6T.M-81)P;1U3e5;?
+R&F\I-Y3\<.WIO7NBZ(DM#Y_[)OL3SOSEQXXWB&P;-X9A5UFQ@,4B3CY<.@#NX?
R&9=X<8E5DT3B,4e0e=JG0&/cIQ\;3_QaO5\(1J_I,(bB\dE^cH[O1L2<0.U<,25
f(#eT:RGD3XH0,GF&DbOF5K9c3GD>9A#2EVL0<9X]EE28>NM@0TS&CQ-GU[W3c5O
;=Y1)N22cLXN,@W\cCHPX[=EA+P[b<X0R(57d.H+\[P7a];@1#<N7B#)-R:Y_4&:
MKBbYE@L1a_4@89DONSM-Ye#<>AJ/-K4)+NX\O:-B(QJZ\fSef@\W2Y+P_&0>Kf7
;dYLgB_:M].]VUI+PKb3R(X.00XeV>&IQ>KD@;g@_?fe-N7/25f]+-^aF3a#a&S7
LK@Od)TE?AFA>Z#:A2)-]Q:.ZK&8g.cHD=3006<D-0EB1&]NCNY9+e/>ZP-(Xf=?
f2D7Y&Ne@LMK0AHLd,H=.Z?K-HeJJ(3b:;CVMgKQF]()R8+[A0cRJc4_eF48H4Q>
?4HLcG/GQ6,fJ[ZN/P-eBBOT(\b:,+3/_;b.=;Dda>YD?832]]2MCEd^CMHCIG<R
8@Oge\4@M1F:(^6OM#]:83cMV6.=MMYWf\6,+6g^X2L4Yfg(E=\Y12PM.CJCa;@O
IAE2W.a0X/bMW&4\H+HX78(Yf1QDb-^:[9HDF2,KXC+^\/92T=[5IQBTaPKH8NR(
CdC?LI?_PC/J2W4+7\E8A?e];9;.;LTgDfc7/#_e(.OWU4dA0=5L(K(C)C8>@25<
YS#/P1<K<AE#6f/99EJ/E0?BR>6/?&/ZWcK6C9J?)cJfQ8J]ZE1c:=?7?,R[W&4O
K>/MDY2fQ@C0IJOQR0c[]=#;57bEU3.Y2H:#305-(:)gN1IP5AEKEA3Eag,CfQ2E
_cMBd#5V4:STe2(><UYD<[QR.6^aA@,OGM85>_>HSg03,AR:[eI^@9L>F24-B+P:
JY8DD;8.V8@#<d?WRU5&2JEd+&U1VLR-[M>JaSD8(?OZXM0<K67+#EE),c@F5T_e
K]P^a[6HO&&fZT9#/R_BL8BS,]Ca54WR3OQOHLU:R3+YccQ^LBN=L;4TWCMH;dZ1
<>>Y/LK)&V>;9Tb#EbOLcI-=HCIaG.:#9SeUZKU:0_((PQRNOb@CffZ^_[YO2D8;
V/V[4HcV>OOHWe>YB0fdgZF(./Y6Kf]F>-YL&K,Ne4;:JHDc19COEDA9>83GX;X_
e553FW3?.8.IY]G4<;+WJ2:<&DUGG@+G_7S(U#@?TgCTRfC\C#_UOQ6=463\P;0M
A;^Y9K_T9=bNGTWR#^+\dBb&P)WH3#CSDQe<Ld.fN8=1T)N-&4AO\=;OSAK=-2@&
=SX&EK&U/G.J5@^\Jc@J?TE2>SJYa168SL5T,2(^V0NJ0gW-K+dN?4eY2612Y=0C
d29?Q2>b-CHDH2N\5B\#07A:KN]1aLS,8@6;)XDbWJ/:;3=/S814VE7]-4C#TN=Q
UJSP\KM^0=GYT5-7^,(TVW_0CU]U>IY<KGSI()?TfX&ZS@gd0CV]Q^0>N1P=+N1M
>)LV4,e[;E..GG:W#YbYB0KN:Z.)+D\g=?aG4&S2a#2QD,CYaH]C-c?4<4)#ST27
2P<SS-N_UQ_::8_dgD<[VYM45beg&>6-R/+/f=6^AZ<6H_dRbYSFg;JOd@ZCVU,@
9UQ0a\;Ke_^?EPF/g/-7?e<[R(-K3;07=@05(Zc&;2>e<[2.IeIf&>gQ(\Z\-KL&
-W+;Q8)c^SEI70_(AbI#9F.60.RD/230E+L#c4(/1_GK_#]f(FQLH:A7>d98MJbR
IMc6cI,EJ)eaQZGMHc/(H[6FZ<+f(4ARCd2I#?CJE\_>=eT9Xg4fE\RV#[g.A4.7
I[Z<J=fg..)X?)+NG#B]^::LVY,LRR+28;N^4=GE)c=E[6[UNWAQ[M9>@VV#J7cI
3DDN3#H>ER/0TNc6BQ-S5J4@=4#=^a0^>4c&1d[SQ?PLMBa5@1]aa9,-:XeM]BY^
,]ULM2&8-BFWZbSY2>KJ^Kf/HW&8e)2dJX>E(1+IE;gA_<\f9fNg).\EUU4@50@]
U.cC@Y1L-[68(Ea/J6K<e/Q0);YReC1X6K\f1GdP<#@-V4@.D=cd]J_(_SG=gTZT
5WEU\DJZ)<XWbT))-^G3-M>]L0W:T4DR2V6.6])P/M@5KdSU)d85]Y&;a.:,_5>F
HRQ2UXX98H_L.6M/dQSN+TIS#X5A^3O[C76aS(be98QdX?JYKGK7cCE.C9@Ib[g\
d+&X^VETSdISE[RN>NPQO#WdT,A(EK0X?F8>4C8?B7/EP-T(:OF\/PN\>J4Kgg@M
&(Od[)UT:P&/>.YR9R2[SYHZe0N,#TB;3#5DG/ZAYR8FBJH.),Z4.PH?]]RNXBTL
KR9\)G0_3(+7Eg#R<?+7+=98)e[(#+O1f;_=8a=_:8QNB:GN/+@eH:#)#^77@P1[
X<Vc:)_,HO=J^-@M],M[R:=TU]X<)1bHCf1I0.KT(]UaP(\6G9&?WbKFW].1(O^=
KXbeCe+8PZ^IT@]JgH#2IO\@b0I+1B<DALIGa?_\[&bE#2bL3.B)-OdU32e8b\a-
P<:5OFIEQ1#6L2Z@&I>X<^RUR^UMA;(YKIP@7A4XM:EQI^fLIABI7.\I<=K3G[H4
37fL;])E,Q\<KgAOJ/:Q1;4(\Ed,[.?JgU9HcDPL;QN:;&X)]bIU\IGU79=4Ve7\
8HTDRXJ^F_J66Be2+2.Y3&?EGO1LJ?1X)\:aU0/C/86,F6-58fI(/RIO_8-dCOGc
3797XTb?FY^F6P)ge+Z>\=c=SPQWZ/<8TY4[.FgW_SVP-E_VaZD0c(F#5/O,N.ge
QW=;9@-FCZ<;SE3D[:K8cSa)6).]W(\dZR,CD4b\3:K49C0Va4,7;e972YOf,^FD
Z<PN7<DU?IZI^>a)590HKVK&.fBPD1LF-IB<7c;2S-M7#-J\M37IWF2>(?^?RW5M
[9b(O)f[a3KUd>7TZ)T6APGCZ62/B(/5TV#T7X3J2T##c;3:KF3Q1JJd-.GIYC(Q
,)].\)6MTF],cb/a?_7CVa<O/&B5DCW9A0=&?a.aLYQ1GEO4R#c3&Q&S;MUK5L=?
\d_F.F^+84@6eRB;CE]V&Z#gV82K=cE5+/YP4\@.bO+XXWZ:.;E@WKLIBBd5PbFK
2bG4NCc[[L2LN7(S>:X+.H6R5I@dGAX\)(KDDfe0B#Z(Tc)E1L,/7)4fTEfBIa0C
1HD^N<&ME.0RfCA)@0aTXVU\02C6M1QM/.FJ/cHQUI?9aP75d0Q+@90]5Lf]8ZQ]
;K?1<>9BgFZ6:(DK\H+:T;D+a=,K[7LRc@N>(H^SHPQeTB^YH<cbY348G/.E4L\T
e_I]IIPg]MNP1575CK9b\\)6DWZI#/GWI.PXM(.&9(J;X1(^K\#:^[+O6J:@KF1L
NQAZf,?W-99>V8e,8JTf?+4J5c(LA,g&EKGE?FYZ57?,.;J@Se1FG:4CTG=()X35
f)TcAI3P7,1]M1/JDC>H,JX)#V.@YHaXH,[eOL-2c^B[d@567I;<XA.AY.DcV_(0
7e[=;FGS2/^Eeg=Xc@6GH[#dCGO-;.Df\O)3^->U0&<,U#V)dIS(f32](g5=<RKT
NK3+\<[;2I>#M.^-^2K0VT37WNb\B8P]H>64^SN4;)>&;0cW9]5bc=>X/FC4b3e@
5S:[JD_MH:9:U?3RA^5=^0EM2KGSe)#0Age5FN;,7XgYXF78I]-)[+fULA[U;+b&
BDOW]6DbG0Z>0e&.g[(XXe1Y_+S-6?>M^(AIU0V\:/D[Ua\0/8-7MUTf24a7[,K^
NVW6-Z>g/YX3MO5S5.<G>88SY0^c>JS^4:NAA5MgN#B#T@.6Y^MYYfYa2Q8CIDG1
4U#<,Y]RKOd<ga#/b_W,,YXOEO]VJ?=aJXda-S)TKD1^^XJIcKSePJ^@_&PbOPPK
c666c;6<[JGDa2L;NI5e-X&[IZ1_df^5GAT/GZT3C.ITA?^^S+XMK_&HPf]8ZYc[
8.Zc[CcR@-^)+WQ^g52@/BG<1U/#^@N_F_G9-Z^/1@0[AHbFIG=LN_N[_TO@FRF/
bc0X=<P/^?]ZbXLC0GE@L(\Mg_.A32:H2DOL]TBcEZ6<7]HP>0Q<>7\1ND\[8?QO
<<B@)\e\D[:@F\/TF9=B-/_f0\=;BAOI)X._ASRJ@fP+4+Z9E:EZ8T[B_)H7:a>&
IF8]MP^g22aJ9(eG/IDEA2]Q>O6LEKRIMJ:Z;U+Oa&W))FDZaC4FdLXd&Cc)gRdY
e63IR)L3<ETK@DT:.NfCN=R&M1Q(60bK<06NK8142E(BK[PZ5Nd&WT/cX<9\M+S=
c;b(#__@(S0&68;F2QBfCL7(:&/.A6UOG^,R(H3I/9dYP[)d.>J:U\-)O:Z.IL-3
9LdUQL)&YXNT5B5SHT2UCA98;M5>&.9C;[D>ZP19^L&+XG5>#(3U,U3LX6G>.G]-
fBO+#K&#[)FD]d-FUMW.\gCB^@]f\2[\+BF/g/D[aE#LeH8SWbHg_21I.8PM7UTb
@;(=(Z94f<TU;[d8W73Xc#41F6V=_eP2Y^6+I77S^C[5e;Q9M?bMV-BK2CY2MdJO
B&)2\&3ec+=da,\:T]3H7gH9K@5Pf,+V<7F8.&39E?&,Idd(-CCWa_X5.97gCHf(
R&F2[TaGJbJP:f.QV?gZ3Tg>DQg<)gW1+c#+3ZILS)fO+(+cY--FWT<4b\e2AS>0
bF;483a0dfg.c9/dI-;BI9EFHVZ81PPD)G0Nd17?G<MAE3G>@_X)Q9O.6dI_1JUc
4E.a&AaI5T)fD(0D)3&A+9gL-@MEB#Nd7NW1,R)T3:&,Z\UYPa@=Mc5AEPM3cHR>
L^[QK[\e4gCg2,O\YD7RgO;ecSK);^-SR/Lg8#&>U,>0KZc[,YcSGC8B:\<8gFY9
K5MIXLd,-YUMWP<E/SgUeWPXYDWF&0e4;W-+LN\]f8[bZAbbC6Q&ZAcG^2Dg^=Fe
MI-[LP[6\B3,1f8ZEFcKTPP6R;0ERAbVZG^<FB^O>>(?_Q8,TO:g</&Q6,Q@UVaJ
:9+=K^ec;;fQ33==J+NLTJ@17Q>e,1c6RB^abIc65X0SaE4J8K6e=HNE]DE#3H0a
5MTgQe=2ac0P]?9Q<RMZ3<^P8Ee3Dga0<D6U,)+.f[..<Xd6:E0/+3+W[,K@6.KW
3KA<#=cXWGQ0<1_9T4O/SbcSHBd4?LS:V64?:FBJ?b2C1D]e@U]gK#Og3<GAWJP(
E.Y@1bQ,\M3+?78@NJ2W8M^91e#3F0=c_RG<0[VSaD@2J8/E#\85IbPbT[@&G>00
O,OVA>e0/-dT\4f0K8Y^OQ.D7?BENSU\f=B6#2_(f2Tf,(5IWN]QSePMD>S@SR6F
/Uf0Z3/dabcO+eCN_G[F3_GVQVd9XODX(+_5LV1BVPOa5GG>cKa(Y:ReXa4;P04F
/Q[JLKR(^ZSCfN<(/T-dFCd+2FFNNNbc=2.9>G&:H(;QMR?1b4<[c5WRNgc9G=+J
DN6#DXVQ)87[,OB[GdE@1-C>AC,8SBb4BEZYWT+RU<MH9ZM18PQLH1c>;KU);5WM
fg<EfW#YdAX(MRKLIKC4#SY29B.3?AE\5_9,UdL(f?c\Q/W<.@NC5(VFAQFRWI[7
OB3VIdJ4[2U3QgC8\-K2XL-@29__@]U/,gG36Y2C-:1b?MfP7#Xb67_OFM<;P\4^
DCF3G1)Z;C>7^@SW7bae:^W?\+S#MNfZ3LL:1=WC)W0B))=H2L>AYOa7L=?W=T.J
#TKMEe(<]7+8>[7BJ\?YLc-/4MH>g:E2NQ;0CL#[@^QH#:b\OD:\CKBWHKJfAO;O
DXK^8V1=T\86H[TJKA9DHK8S//eH\G<W43df=Wg;SH3gVBb=a>-?cg=.Zc;YSSF@
_LD0EM+>)Ue6AKCMVP><ZbCH_6XKRPY,@[R)dDH,,F5U-]P7O+16c&)7>499A2b4
>\QD.1^LbW>DZ/?[CPCJUXF7C<R>5]PFW)50N44cYa.-G,EUUZ?/11^N6>WK;aW2
PELU8Q4[I@bRW(#);ZTgZgaYe+\/?\?;#0IU.CLZYL.7N://-5P)&UJOSg2+LA)e
LE3a=b7;.?a9CIQ[MD+&RU7-[T=CWW-;4a;AOEM<]TTDdDL2:;[_)@8MLHU;2IFf
&\)QaG^Y5Gc-Ge?I8F(XedU?YO1c/)3PP@9G95UP?:C<BV:^OFZ.F\-C6>VS^E)&
5[&R/@IAc::H+CWL^5[3@Qd8&Qaa([[R^8e@3-9A6JN.,bLJ+40@4C+>B-=58aR&
-K4TP,?BDMSV@-6/b[O/AJK&VJYL49+L\cEI(FZ=DTP.+GQYZ,_9fgL)5_91>eVV
3SM3<[0FK5b,JSgG<&.QP9_<T7/a3(gO/_dRDV@YJJ#bQ./7S7e0B<RX1a_1S1C;
1HQNB]<A+&fde[1PT0H^;N9?G[cE1QF/HWE_A/?FW?S7BBcgX:_GB:I\KWR#2Qa)
?G.fU==G^=X#USP6eM.LD[M[]RVZ-575+__6.JWLc?6[O2HN+607DUgc:((^+GGV
L#NBV^ESW3PcBf-f:cKC8)2<LJ5&:V3F&ZC7NOF.TUVI@X^4NTP7<bW=AH,daf-9
IA+1-3ZXV/J^IJQ1d?-\>?KS1B<\N\Z]IRT[6c^)(R-6;OK(0aL,N5^:D_a<;+P)
b]JeJXOBTH<OH9fBT=bVEJ@3?L..bF_@;$
`endprotected


